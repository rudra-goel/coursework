* SPICE NETLIST
***************************************

.SUBCKT 16_bit_ripple_carry_adder gnd! B<1> B<3> B<5> B<7> A<0> A<2> A<4> A<6> A<1> A<3> A<5> A<7> B<0> B<2> B<4> B<6> Sout<1> Sout<3> Sout<5>
+ Sout<7> Sout<0> Sout<2> Sout<4> Sout<6> Cin vdd! B<9> B<11> B<13> B<15> A<8> A<10> A<12> A<14> A<9> A<11> A<13> A<15> B<8>
+ B<10> B<12> B<14> Sout<9> Sout<11> Sout<13> Sout<15> Sout<8> Sout<10> Sout<12> Sout<14> Cout
** N=355 EP=52 IP=0 FDC=576
M0 276 B<1> 6 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=8.82e-14 AS=8.595e-14 PD=1.34e-06 PS=1.315e-06 $X=1530 $Y=6675 $D=1
M1 277 B<3> 7 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=8.82e-14 AS=8.595e-14 PD=1.34e-06 PS=1.315e-06 $X=1530 $Y=14075 $D=1
M2 278 B<5> 8 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=8.82e-14 AS=8.595e-14 PD=1.34e-06 PS=1.315e-06 $X=1530 $Y=21475 $D=1
M3 279 B<7> 9 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=8.82e-14 AS=8.595e-14 PD=1.34e-06 PS=1.315e-06 $X=1530 $Y=28875 $D=1
M4 131 A<0> gnd! gnd! NMOS_VTL L=5e-08 W=9e-08 AD=5.175e-14 AS=5.175e-14 PD=1.33e-06 PS=1.33e-06 $X=1950 $Y=790 $D=1
M5 132 A<2> gnd! gnd! NMOS_VTL L=5e-08 W=9e-08 AD=5.175e-14 AS=5.175e-14 PD=1.33e-06 PS=1.33e-06 $X=1950 $Y=8190 $D=1
M6 133 A<4> gnd! gnd! NMOS_VTL L=5e-08 W=9e-08 AD=5.175e-14 AS=5.175e-14 PD=1.33e-06 PS=1.33e-06 $X=1950 $Y=15590 $D=1
M7 134 A<6> gnd! gnd! NMOS_VTL L=5e-08 W=9e-08 AD=5.175e-14 AS=5.175e-14 PD=1.33e-06 PS=1.33e-06 $X=1950 $Y=22990 $D=1
M8 gnd! A<1> 276 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=7.155e-14 AS=8.82e-14 PD=1.155e-06 PS=1.34e-06 $X=2610 $Y=6675 $D=1
M9 gnd! A<3> 277 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=7.155e-14 AS=8.82e-14 PD=1.155e-06 PS=1.34e-06 $X=2610 $Y=14075 $D=1
M10 gnd! A<5> 278 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=7.155e-14 AS=8.82e-14 PD=1.155e-06 PS=1.34e-06 $X=2610 $Y=21475 $D=1
M11 gnd! A<7> 279 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=7.155e-14 AS=8.82e-14 PD=1.155e-06 PS=1.34e-06 $X=2610 $Y=28875 $D=1
M12 gnd! A<0> 22 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.2285e-13 AS=4.05e-14 PD=1.725e-06 PS=8.1e-07 $X=5350 $Y=900 $D=1
M13 gnd! A<2> 23 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.2285e-13 AS=4.05e-14 PD=1.725e-06 PS=8.1e-07 $X=5350 $Y=8300 $D=1
M14 gnd! A<4> 24 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.2285e-13 AS=4.05e-14 PD=1.725e-06 PS=8.1e-07 $X=5350 $Y=15700 $D=1
M15 gnd! A<6> 25 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.2285e-13 AS=4.05e-14 PD=1.725e-06 PS=8.1e-07 $X=5350 $Y=23100 $D=1
M16 280 6 20 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=8.82e-14 AS=8.595e-14 PD=1.34e-06 PS=1.315e-06 $X=5530 $Y=6675 $D=1
M17 281 7 18 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=8.82e-14 AS=8.595e-14 PD=1.34e-06 PS=1.315e-06 $X=5530 $Y=14075 $D=1
M18 282 8 21 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=8.82e-14 AS=8.595e-14 PD=1.34e-06 PS=1.315e-06 $X=5530 $Y=21475 $D=1
M19 283 9 19 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=8.82e-14 AS=8.595e-14 PD=1.34e-06 PS=1.315e-06 $X=5530 $Y=28875 $D=1
M20 gnd! 135 280 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=7.155e-14 AS=8.82e-14 PD=1.155e-06 PS=1.34e-06 $X=6610 $Y=6675 $D=1
M21 gnd! 136 281 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=7.155e-14 AS=8.82e-14 PD=1.155e-06 PS=1.34e-06 $X=6610 $Y=14075 $D=1
M22 gnd! 137 282 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=7.155e-14 AS=8.82e-14 PD=1.155e-06 PS=1.34e-06 $X=6610 $Y=21475 $D=1
M23 gnd! 138 283 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=7.155e-14 AS=8.82e-14 PD=1.155e-06 PS=1.34e-06 $X=6610 $Y=28875 $D=1
M24 284 143 gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=9.855e-14 AS=1.2285e-13 PD=1.455e-06 PS=1.725e-06 $X=6815 $Y=900 $D=1
M25 285 144 gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=9.855e-14 AS=1.2285e-13 PD=1.455e-06 PS=1.725e-06 $X=6815 $Y=8300 $D=1
M26 286 145 gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=9.855e-14 AS=1.2285e-13 PD=1.455e-06 PS=1.725e-06 $X=6815 $Y=15700 $D=1
M27 287 146 gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=9.855e-14 AS=1.2285e-13 PD=1.455e-06 PS=1.725e-06 $X=6815 $Y=23100 $D=1
M28 26 131 284 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.161e-13 AS=9.855e-14 PD=1.65e-06 PS=1.455e-06 $X=8010 $Y=900 $D=1
M29 27 132 285 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.161e-13 AS=9.855e-14 PD=1.65e-06 PS=1.455e-06 $X=8010 $Y=8300 $D=1
M30 28 133 286 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.161e-13 AS=9.855e-14 PD=1.65e-06 PS=1.455e-06 $X=8010 $Y=15700 $D=1
M31 29 134 287 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.161e-13 AS=9.855e-14 PD=1.65e-06 PS=1.455e-06 $X=8010 $Y=23100 $D=1
M32 22 B<0> 26 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.26e-13 AS=1.161e-13 PD=1.76e-06 PS=1.65e-06 $X=9400 $Y=900 $D=1
M33 23 B<2> 27 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.26e-13 AS=1.161e-13 PD=1.76e-06 PS=1.65e-06 $X=9400 $Y=8300 $D=1
M34 24 B<4> 28 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.26e-13 AS=1.161e-13 PD=1.76e-06 PS=1.65e-06 $X=9400 $Y=15700 $D=1
M35 25 B<6> 29 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.26e-13 AS=1.161e-13 PD=1.76e-06 PS=1.65e-06 $X=9400 $Y=23100 $D=1
M36 288 30 135 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=8.82e-14 AS=8.595e-14 PD=1.34e-06 PS=1.315e-06 $X=9530 $Y=6675 $D=1
M37 289 31 136 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=8.82e-14 AS=8.595e-14 PD=1.34e-06 PS=1.315e-06 $X=9530 $Y=14075 $D=1
M38 290 32 137 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=8.82e-14 AS=8.595e-14 PD=1.34e-06 PS=1.315e-06 $X=9530 $Y=21475 $D=1
M39 291 33 138 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=8.82e-14 AS=8.595e-14 PD=1.34e-06 PS=1.315e-06 $X=9530 $Y=28875 $D=1
M40 gnd! 34 288 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=7.155e-14 AS=8.82e-14 PD=1.155e-06 PS=1.34e-06 $X=10610 $Y=6675 $D=1
M41 gnd! 35 289 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=7.155e-14 AS=8.82e-14 PD=1.155e-06 PS=1.34e-06 $X=10610 $Y=14075 $D=1
M42 gnd! 36 290 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=7.155e-14 AS=8.82e-14 PD=1.155e-06 PS=1.34e-06 $X=10610 $Y=21475 $D=1
M43 gnd! 37 291 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=7.155e-14 AS=8.82e-14 PD=1.155e-06 PS=1.34e-06 $X=10610 $Y=28875 $D=1
M44 gnd! 30 139 gnd! NMOS_VTL L=5e-08 W=9e-08 AD=5.175e-14 AS=5.175e-14 PD=1.33e-06 PS=1.33e-06 $X=13835 $Y=6755 $D=1
M45 gnd! 31 140 gnd! NMOS_VTL L=5e-08 W=9e-08 AD=5.175e-14 AS=5.175e-14 PD=1.33e-06 PS=1.33e-06 $X=13835 $Y=14155 $D=1
M46 gnd! 32 141 gnd! NMOS_VTL L=5e-08 W=9e-08 AD=5.175e-14 AS=5.175e-14 PD=1.33e-06 PS=1.33e-06 $X=13835 $Y=21555 $D=1
M47 gnd! 33 142 gnd! NMOS_VTL L=5e-08 W=9e-08 AD=5.175e-14 AS=5.175e-14 PD=1.33e-06 PS=1.33e-06 $X=13835 $Y=28955 $D=1
M48 143 B<0> gnd! gnd! NMOS_VTL L=5e-08 W=9e-08 AD=5.175e-14 AS=5.175e-14 PD=1.33e-06 PS=1.33e-06 $X=14565 $Y=795 $D=1
M49 144 B<2> gnd! gnd! NMOS_VTL L=5e-08 W=9e-08 AD=5.175e-14 AS=5.175e-14 PD=1.33e-06 PS=1.33e-06 $X=14565 $Y=8195 $D=1
M50 145 B<4> gnd! gnd! NMOS_VTL L=5e-08 W=9e-08 AD=5.175e-14 AS=5.175e-14 PD=1.33e-06 PS=1.33e-06 $X=14565 $Y=15595 $D=1
M51 146 B<6> gnd! gnd! NMOS_VTL L=5e-08 W=9e-08 AD=5.175e-14 AS=5.175e-14 PD=1.33e-06 PS=1.33e-06 $X=14565 $Y=22995 $D=1
M52 147 26 gnd! gnd! NMOS_VTL L=5e-08 W=9e-08 AD=5.175e-14 AS=5.175e-14 PD=1.33e-06 PS=1.33e-06 $X=18450 $Y=790 $D=1
M53 148 27 gnd! gnd! NMOS_VTL L=5e-08 W=9e-08 AD=5.175e-14 AS=5.175e-14 PD=1.33e-06 PS=1.33e-06 $X=18450 $Y=8190 $D=1
M54 149 28 gnd! gnd! NMOS_VTL L=5e-08 W=9e-08 AD=5.175e-14 AS=5.175e-14 PD=1.33e-06 PS=1.33e-06 $X=18450 $Y=15590 $D=1
M55 150 29 gnd! gnd! NMOS_VTL L=5e-08 W=9e-08 AD=5.175e-14 AS=5.175e-14 PD=1.33e-06 PS=1.33e-06 $X=18450 $Y=22990 $D=1
M56 Sout<1> 30 42 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.161e-13 AS=1.26e-13 PD=1.65e-06 PS=1.76e-06 $X=19000 $Y=6470 $D=1
M57 Sout<3> 31 43 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.161e-13 AS=1.26e-13 PD=1.65e-06 PS=1.76e-06 $X=19000 $Y=13870 $D=1
M58 Sout<5> 32 44 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.161e-13 AS=1.26e-13 PD=1.65e-06 PS=1.76e-06 $X=19000 $Y=21270 $D=1
M59 Sout<7> 33 45 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.161e-13 AS=1.26e-13 PD=1.65e-06 PS=1.76e-06 $X=19000 $Y=28670 $D=1
M60 292 151 Sout<1> gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=9.855e-14 AS=1.161e-13 PD=1.455e-06 PS=1.65e-06 $X=20390 $Y=6470 $D=1
M61 293 152 Sout<3> gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=9.855e-14 AS=1.161e-13 PD=1.455e-06 PS=1.65e-06 $X=20390 $Y=13870 $D=1
M62 294 153 Sout<5> gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=9.855e-14 AS=1.161e-13 PD=1.455e-06 PS=1.65e-06 $X=20390 $Y=21270 $D=1
M63 295 154 Sout<7> gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=9.855e-14 AS=1.161e-13 PD=1.455e-06 PS=1.65e-06 $X=20390 $Y=28670 $D=1
M64 gnd! 139 292 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.2285e-13 AS=9.855e-14 PD=1.725e-06 PS=1.455e-06 $X=21585 $Y=6470 $D=1
M65 gnd! 140 293 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.2285e-13 AS=9.855e-14 PD=1.725e-06 PS=1.455e-06 $X=21585 $Y=13870 $D=1
M66 gnd! 141 294 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.2285e-13 AS=9.855e-14 PD=1.725e-06 PS=1.455e-06 $X=21585 $Y=21270 $D=1
M67 gnd! 142 295 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.2285e-13 AS=9.855e-14 PD=1.725e-06 PS=1.455e-06 $X=21585 $Y=28670 $D=1
M68 gnd! 26 50 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.2285e-13 AS=4.05e-14 PD=1.725e-06 PS=8.1e-07 $X=21850 $Y=900 $D=1
M69 gnd! 27 51 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.2285e-13 AS=4.05e-14 PD=1.725e-06 PS=8.1e-07 $X=21850 $Y=8300 $D=1
M70 gnd! 28 52 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.2285e-13 AS=4.05e-14 PD=1.725e-06 PS=8.1e-07 $X=21850 $Y=15700 $D=1
M71 gnd! 29 53 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.2285e-13 AS=4.05e-14 PD=1.725e-06 PS=8.1e-07 $X=21850 $Y=23100 $D=1
M72 42 34 gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=4.05e-14 AS=1.2285e-13 PD=8.1e-07 PS=1.725e-06 $X=23050 $Y=6470 $D=1
M73 43 35 gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=4.05e-14 AS=1.2285e-13 PD=8.1e-07 PS=1.725e-06 $X=23050 $Y=13870 $D=1
M74 44 36 gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=4.05e-14 AS=1.2285e-13 PD=8.1e-07 PS=1.725e-06 $X=23050 $Y=21270 $D=1
M75 45 37 gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=4.05e-14 AS=1.2285e-13 PD=8.1e-07 PS=1.725e-06 $X=23050 $Y=28670 $D=1
M76 296 159 gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=9.855e-14 AS=1.2285e-13 PD=1.455e-06 PS=1.725e-06 $X=23315 $Y=900 $D=1
M77 297 160 gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=9.855e-14 AS=1.2285e-13 PD=1.455e-06 PS=1.725e-06 $X=23315 $Y=8300 $D=1
M78 298 161 gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=9.855e-14 AS=1.2285e-13 PD=1.455e-06 PS=1.725e-06 $X=23315 $Y=15700 $D=1
M79 299 162 gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=9.855e-14 AS=1.2285e-13 PD=1.455e-06 PS=1.725e-06 $X=23315 $Y=23100 $D=1
M80 Sout<0> 147 296 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.161e-13 AS=9.855e-14 PD=1.65e-06 PS=1.455e-06 $X=24510 $Y=900 $D=1
M81 Sout<2> 148 297 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.161e-13 AS=9.855e-14 PD=1.65e-06 PS=1.455e-06 $X=24510 $Y=8300 $D=1
M82 Sout<4> 149 298 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.161e-13 AS=9.855e-14 PD=1.65e-06 PS=1.455e-06 $X=24510 $Y=15700 $D=1
M83 Sout<6> 150 299 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.161e-13 AS=9.855e-14 PD=1.65e-06 PS=1.455e-06 $X=24510 $Y=23100 $D=1
M84 50 Cin Sout<0> gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.26e-13 AS=1.161e-13 PD=1.76e-06 PS=1.65e-06 $X=25900 $Y=900 $D=1
M85 51 20 Sout<2> gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.26e-13 AS=1.161e-13 PD=1.76e-06 PS=1.65e-06 $X=25900 $Y=8300 $D=1
M86 52 18 Sout<4> gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.26e-13 AS=1.161e-13 PD=1.76e-06 PS=1.65e-06 $X=25900 $Y=15700 $D=1
M87 53 21 Sout<6> gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.26e-13 AS=1.161e-13 PD=1.76e-06 PS=1.65e-06 $X=25900 $Y=23100 $D=1
M88 gnd! 34 151 gnd! NMOS_VTL L=5e-08 W=9e-08 AD=5.175e-14 AS=5.175e-14 PD=1.33e-06 PS=1.33e-06 $X=26450 $Y=6760 $D=1
M89 gnd! 35 152 gnd! NMOS_VTL L=5e-08 W=9e-08 AD=5.175e-14 AS=5.175e-14 PD=1.33e-06 PS=1.33e-06 $X=26450 $Y=14160 $D=1
M90 gnd! 36 153 gnd! NMOS_VTL L=5e-08 W=9e-08 AD=5.175e-14 AS=5.175e-14 PD=1.33e-06 PS=1.33e-06 $X=26450 $Y=21560 $D=1
M91 gnd! 37 154 gnd! NMOS_VTL L=5e-08 W=9e-08 AD=5.175e-14 AS=5.175e-14 PD=1.33e-06 PS=1.33e-06 $X=26450 $Y=28960 $D=1
M92 gnd! B<1> 155 gnd! NMOS_VTL L=5e-08 W=9e-08 AD=5.175e-14 AS=5.175e-14 PD=1.33e-06 PS=1.33e-06 $X=30335 $Y=6755 $D=1
M93 gnd! B<3> 156 gnd! NMOS_VTL L=5e-08 W=9e-08 AD=5.175e-14 AS=5.175e-14 PD=1.33e-06 PS=1.33e-06 $X=30335 $Y=14155 $D=1
M94 gnd! B<5> 157 gnd! NMOS_VTL L=5e-08 W=9e-08 AD=5.175e-14 AS=5.175e-14 PD=1.33e-06 PS=1.33e-06 $X=30335 $Y=21555 $D=1
M95 gnd! B<7> 158 gnd! NMOS_VTL L=5e-08 W=9e-08 AD=5.175e-14 AS=5.175e-14 PD=1.33e-06 PS=1.33e-06 $X=30335 $Y=28955 $D=1
M96 159 Cin gnd! gnd! NMOS_VTL L=5e-08 W=9e-08 AD=5.175e-14 AS=5.175e-14 PD=1.33e-06 PS=1.33e-06 $X=31065 $Y=795 $D=1
M97 160 20 gnd! gnd! NMOS_VTL L=5e-08 W=9e-08 AD=5.175e-14 AS=5.175e-14 PD=1.33e-06 PS=1.33e-06 $X=31065 $Y=8195 $D=1
M98 161 18 gnd! gnd! NMOS_VTL L=5e-08 W=9e-08 AD=5.175e-14 AS=5.175e-14 PD=1.33e-06 PS=1.33e-06 $X=31065 $Y=15595 $D=1
M99 162 21 gnd! gnd! NMOS_VTL L=5e-08 W=9e-08 AD=5.175e-14 AS=5.175e-14 PD=1.33e-06 PS=1.33e-06 $X=31065 $Y=22995 $D=1
M100 300 26 gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=8.82e-14 AS=7.155e-14 PD=1.34e-06 PS=1.155e-06 $X=34290 $Y=695 $D=1
M101 301 27 gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=8.82e-14 AS=7.155e-14 PD=1.34e-06 PS=1.155e-06 $X=34290 $Y=8095 $D=1
M102 302 28 gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=8.82e-14 AS=7.155e-14 PD=1.34e-06 PS=1.155e-06 $X=34290 $Y=15495 $D=1
M103 303 29 gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=8.82e-14 AS=7.155e-14 PD=1.34e-06 PS=1.155e-06 $X=34290 $Y=22895 $D=1
M104 163 Cin 300 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=8.595e-14 AS=8.82e-14 PD=1.315e-06 PS=1.34e-06 $X=35370 $Y=695 $D=1
M105 164 20 301 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=8.595e-14 AS=8.82e-14 PD=1.315e-06 PS=1.34e-06 $X=35370 $Y=8095 $D=1
M106 165 18 302 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=8.595e-14 AS=8.82e-14 PD=1.315e-06 PS=1.34e-06 $X=35370 $Y=15495 $D=1
M107 166 21 303 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=8.595e-14 AS=8.82e-14 PD=1.315e-06 PS=1.34e-06 $X=35370 $Y=22895 $D=1
M108 34 B<1> 59 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.161e-13 AS=1.26e-13 PD=1.65e-06 PS=1.76e-06 $X=35500 $Y=6470 $D=1
M109 35 B<3> 60 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.161e-13 AS=1.26e-13 PD=1.65e-06 PS=1.76e-06 $X=35500 $Y=13870 $D=1
M110 36 B<5> 61 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.161e-13 AS=1.26e-13 PD=1.65e-06 PS=1.76e-06 $X=35500 $Y=21270 $D=1
M111 37 B<7> 62 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.161e-13 AS=1.26e-13 PD=1.65e-06 PS=1.76e-06 $X=35500 $Y=28670 $D=1
M112 304 167 34 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=9.855e-14 AS=1.161e-13 PD=1.455e-06 PS=1.65e-06 $X=36890 $Y=6470 $D=1
M113 305 168 35 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=9.855e-14 AS=1.161e-13 PD=1.455e-06 PS=1.65e-06 $X=36890 $Y=13870 $D=1
M114 306 169 36 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=9.855e-14 AS=1.161e-13 PD=1.455e-06 PS=1.65e-06 $X=36890 $Y=21270 $D=1
M115 307 170 37 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=9.855e-14 AS=1.161e-13 PD=1.455e-06 PS=1.65e-06 $X=36890 $Y=28670 $D=1
M116 gnd! 155 304 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.2285e-13 AS=9.855e-14 PD=1.725e-06 PS=1.455e-06 $X=38085 $Y=6470 $D=1
M117 gnd! 156 305 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.2285e-13 AS=9.855e-14 PD=1.725e-06 PS=1.455e-06 $X=38085 $Y=13870 $D=1
M118 gnd! 157 306 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.2285e-13 AS=9.855e-14 PD=1.725e-06 PS=1.455e-06 $X=38085 $Y=21270 $D=1
M119 gnd! 158 307 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.2285e-13 AS=9.855e-14 PD=1.725e-06 PS=1.455e-06 $X=38085 $Y=28670 $D=1
M120 308 163 gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=8.82e-14 AS=7.155e-14 PD=1.34e-06 PS=1.155e-06 $X=38290 $Y=695 $D=1
M121 309 164 gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=8.82e-14 AS=7.155e-14 PD=1.34e-06 PS=1.155e-06 $X=38290 $Y=8095 $D=1
M122 310 165 gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=8.82e-14 AS=7.155e-14 PD=1.34e-06 PS=1.155e-06 $X=38290 $Y=15495 $D=1
M123 311 166 gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=8.82e-14 AS=7.155e-14 PD=1.34e-06 PS=1.155e-06 $X=38290 $Y=22895 $D=1
M124 30 63 308 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=8.595e-14 AS=8.82e-14 PD=1.315e-06 PS=1.34e-06 $X=39370 $Y=695 $D=1
M125 31 64 309 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=8.595e-14 AS=8.82e-14 PD=1.315e-06 PS=1.34e-06 $X=39370 $Y=8095 $D=1
M126 32 65 310 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=8.595e-14 AS=8.82e-14 PD=1.315e-06 PS=1.34e-06 $X=39370 $Y=15495 $D=1
M127 33 66 311 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=8.595e-14 AS=8.82e-14 PD=1.315e-06 PS=1.34e-06 $X=39370 $Y=22895 $D=1
M128 59 A<1> gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=4.05e-14 AS=1.2285e-13 PD=8.1e-07 PS=1.725e-06 $X=39550 $Y=6470 $D=1
M129 60 A<3> gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=4.05e-14 AS=1.2285e-13 PD=8.1e-07 PS=1.725e-06 $X=39550 $Y=13870 $D=1
M130 61 A<5> gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=4.05e-14 AS=1.2285e-13 PD=8.1e-07 PS=1.725e-06 $X=39550 $Y=21270 $D=1
M131 62 A<7> gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=4.05e-14 AS=1.2285e-13 PD=8.1e-07 PS=1.725e-06 $X=39550 $Y=28670 $D=1
M132 312 A<0> gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=8.82e-14 AS=7.155e-14 PD=1.34e-06 PS=1.155e-06 $X=42290 $Y=695 $D=1
M133 313 A<2> gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=8.82e-14 AS=7.155e-14 PD=1.34e-06 PS=1.155e-06 $X=42290 $Y=8095 $D=1
M134 314 A<4> gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=8.82e-14 AS=7.155e-14 PD=1.34e-06 PS=1.155e-06 $X=42290 $Y=15495 $D=1
M135 315 A<6> gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=8.82e-14 AS=7.155e-14 PD=1.34e-06 PS=1.155e-06 $X=42290 $Y=22895 $D=1
M136 gnd! A<1> 167 gnd! NMOS_VTL L=5e-08 W=9e-08 AD=5.175e-14 AS=5.175e-14 PD=1.33e-06 PS=1.33e-06 $X=42950 $Y=6760 $D=1
M137 gnd! A<3> 168 gnd! NMOS_VTL L=5e-08 W=9e-08 AD=5.175e-14 AS=5.175e-14 PD=1.33e-06 PS=1.33e-06 $X=42950 $Y=14160 $D=1
M138 gnd! A<5> 169 gnd! NMOS_VTL L=5e-08 W=9e-08 AD=5.175e-14 AS=5.175e-14 PD=1.33e-06 PS=1.33e-06 $X=42950 $Y=21560 $D=1
M139 gnd! A<7> 170 gnd! NMOS_VTL L=5e-08 W=9e-08 AD=5.175e-14 AS=5.175e-14 PD=1.33e-06 PS=1.33e-06 $X=42950 $Y=28960 $D=1
M140 63 B<0> 312 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=8.595e-14 AS=8.82e-14 PD=1.315e-06 PS=1.34e-06 $X=43370 $Y=695 $D=1
M141 64 B<2> 313 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=8.595e-14 AS=8.82e-14 PD=1.315e-06 PS=1.34e-06 $X=43370 $Y=8095 $D=1
M142 65 B<4> 314 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=8.595e-14 AS=8.82e-14 PD=1.315e-06 PS=1.34e-06 $X=43370 $Y=15495 $D=1
M143 66 B<6> 315 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=8.595e-14 AS=8.82e-14 PD=1.315e-06 PS=1.34e-06 $X=43370 $Y=22895 $D=1
M144 316 B<9> 72 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=8.82e-14 AS=8.595e-14 PD=1.34e-06 PS=1.315e-06 $X=46530 $Y=6675 $D=1
M145 317 B<11> 73 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=8.82e-14 AS=8.595e-14 PD=1.34e-06 PS=1.315e-06 $X=46530 $Y=14075 $D=1
M146 318 B<13> 74 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=8.82e-14 AS=8.595e-14 PD=1.34e-06 PS=1.315e-06 $X=46530 $Y=21475 $D=1
M147 319 B<15> 75 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=8.82e-14 AS=8.595e-14 PD=1.34e-06 PS=1.315e-06 $X=46530 $Y=28875 $D=1
M148 171 A<8> gnd! gnd! NMOS_VTL L=5e-08 W=9e-08 AD=5.175e-14 AS=5.175e-14 PD=1.33e-06 PS=1.33e-06 $X=46950 $Y=790 $D=1
M149 172 A<10> gnd! gnd! NMOS_VTL L=5e-08 W=9e-08 AD=5.175e-14 AS=5.175e-14 PD=1.33e-06 PS=1.33e-06 $X=46950 $Y=8190 $D=1
M150 173 A<12> gnd! gnd! NMOS_VTL L=5e-08 W=9e-08 AD=5.175e-14 AS=5.175e-14 PD=1.33e-06 PS=1.33e-06 $X=46950 $Y=15590 $D=1
M151 174 A<14> gnd! gnd! NMOS_VTL L=5e-08 W=9e-08 AD=5.175e-14 AS=5.175e-14 PD=1.33e-06 PS=1.33e-06 $X=46950 $Y=22990 $D=1
M152 gnd! A<9> 316 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=7.155e-14 AS=8.82e-14 PD=1.155e-06 PS=1.34e-06 $X=47610 $Y=6675 $D=1
M153 gnd! A<11> 317 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=7.155e-14 AS=8.82e-14 PD=1.155e-06 PS=1.34e-06 $X=47610 $Y=14075 $D=1
M154 gnd! A<13> 318 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=7.155e-14 AS=8.82e-14 PD=1.155e-06 PS=1.34e-06 $X=47610 $Y=21475 $D=1
M155 gnd! A<15> 319 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=7.155e-14 AS=8.82e-14 PD=1.155e-06 PS=1.34e-06 $X=47610 $Y=28875 $D=1
M156 gnd! A<8> 87 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.2285e-13 AS=4.05e-14 PD=1.725e-06 PS=8.1e-07 $X=50350 $Y=900 $D=1
M157 gnd! A<10> 88 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.2285e-13 AS=4.05e-14 PD=1.725e-06 PS=8.1e-07 $X=50350 $Y=8300 $D=1
M158 gnd! A<12> 89 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.2285e-13 AS=4.05e-14 PD=1.725e-06 PS=8.1e-07 $X=50350 $Y=15700 $D=1
M159 gnd! A<14> 90 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.2285e-13 AS=4.05e-14 PD=1.725e-06 PS=8.1e-07 $X=50350 $Y=23100 $D=1
M160 320 72 85 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=8.82e-14 AS=8.595e-14 PD=1.34e-06 PS=1.315e-06 $X=50530 $Y=6675 $D=1
M161 321 73 84 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=8.82e-14 AS=8.595e-14 PD=1.34e-06 PS=1.315e-06 $X=50530 $Y=14075 $D=1
M162 322 74 86 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=8.82e-14 AS=8.595e-14 PD=1.34e-06 PS=1.315e-06 $X=50530 $Y=21475 $D=1
M163 323 75 Cout gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=8.82e-14 AS=8.595e-14 PD=1.34e-06 PS=1.315e-06 $X=50530 $Y=28875 $D=1
M164 gnd! 176 320 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=7.155e-14 AS=8.82e-14 PD=1.155e-06 PS=1.34e-06 $X=51610 $Y=6675 $D=1
M165 gnd! 177 321 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=7.155e-14 AS=8.82e-14 PD=1.155e-06 PS=1.34e-06 $X=51610 $Y=14075 $D=1
M166 gnd! 178 322 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=7.155e-14 AS=8.82e-14 PD=1.155e-06 PS=1.34e-06 $X=51610 $Y=21475 $D=1
M167 gnd! 179 323 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=7.155e-14 AS=8.82e-14 PD=1.155e-06 PS=1.34e-06 $X=51610 $Y=28875 $D=1
M168 324 184 gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=9.855e-14 AS=1.2285e-13 PD=1.455e-06 PS=1.725e-06 $X=51815 $Y=900 $D=1
M169 325 185 gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=9.855e-14 AS=1.2285e-13 PD=1.455e-06 PS=1.725e-06 $X=51815 $Y=8300 $D=1
M170 326 186 gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=9.855e-14 AS=1.2285e-13 PD=1.455e-06 PS=1.725e-06 $X=51815 $Y=15700 $D=1
M171 327 187 gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=9.855e-14 AS=1.2285e-13 PD=1.455e-06 PS=1.725e-06 $X=51815 $Y=23100 $D=1
M172 91 171 324 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.161e-13 AS=9.855e-14 PD=1.65e-06 PS=1.455e-06 $X=53010 $Y=900 $D=1
M173 92 172 325 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.161e-13 AS=9.855e-14 PD=1.65e-06 PS=1.455e-06 $X=53010 $Y=8300 $D=1
M174 93 173 326 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.161e-13 AS=9.855e-14 PD=1.65e-06 PS=1.455e-06 $X=53010 $Y=15700 $D=1
M175 94 174 327 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.161e-13 AS=9.855e-14 PD=1.65e-06 PS=1.455e-06 $X=53010 $Y=23100 $D=1
M176 87 B<8> 91 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.26e-13 AS=1.161e-13 PD=1.76e-06 PS=1.65e-06 $X=54400 $Y=900 $D=1
M177 88 B<10> 92 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.26e-13 AS=1.161e-13 PD=1.76e-06 PS=1.65e-06 $X=54400 $Y=8300 $D=1
M178 89 B<12> 93 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.26e-13 AS=1.161e-13 PD=1.76e-06 PS=1.65e-06 $X=54400 $Y=15700 $D=1
M179 90 B<14> 94 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.26e-13 AS=1.161e-13 PD=1.76e-06 PS=1.65e-06 $X=54400 $Y=23100 $D=1
M180 328 95 176 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=8.82e-14 AS=8.595e-14 PD=1.34e-06 PS=1.315e-06 $X=54530 $Y=6675 $D=1
M181 329 96 177 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=8.82e-14 AS=8.595e-14 PD=1.34e-06 PS=1.315e-06 $X=54530 $Y=14075 $D=1
M182 330 97 178 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=8.82e-14 AS=8.595e-14 PD=1.34e-06 PS=1.315e-06 $X=54530 $Y=21475 $D=1
M183 331 98 179 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=8.82e-14 AS=8.595e-14 PD=1.34e-06 PS=1.315e-06 $X=54530 $Y=28875 $D=1
M184 gnd! 99 328 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=7.155e-14 AS=8.82e-14 PD=1.155e-06 PS=1.34e-06 $X=55610 $Y=6675 $D=1
M185 gnd! 100 329 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=7.155e-14 AS=8.82e-14 PD=1.155e-06 PS=1.34e-06 $X=55610 $Y=14075 $D=1
M186 gnd! 101 330 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=7.155e-14 AS=8.82e-14 PD=1.155e-06 PS=1.34e-06 $X=55610 $Y=21475 $D=1
M187 gnd! 102 331 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=7.155e-14 AS=8.82e-14 PD=1.155e-06 PS=1.34e-06 $X=55610 $Y=28875 $D=1
M188 gnd! 95 180 gnd! NMOS_VTL L=5e-08 W=9e-08 AD=5.175e-14 AS=5.175e-14 PD=1.33e-06 PS=1.33e-06 $X=58835 $Y=6755 $D=1
M189 gnd! 96 181 gnd! NMOS_VTL L=5e-08 W=9e-08 AD=5.175e-14 AS=5.175e-14 PD=1.33e-06 PS=1.33e-06 $X=58835 $Y=14155 $D=1
M190 gnd! 97 182 gnd! NMOS_VTL L=5e-08 W=9e-08 AD=5.175e-14 AS=5.175e-14 PD=1.33e-06 PS=1.33e-06 $X=58835 $Y=21555 $D=1
M191 gnd! 98 183 gnd! NMOS_VTL L=5e-08 W=9e-08 AD=5.175e-14 AS=5.175e-14 PD=1.33e-06 PS=1.33e-06 $X=58835 $Y=28955 $D=1
M192 184 B<8> gnd! gnd! NMOS_VTL L=5e-08 W=9e-08 AD=5.175e-14 AS=5.175e-14 PD=1.33e-06 PS=1.33e-06 $X=59565 $Y=795 $D=1
M193 185 B<10> gnd! gnd! NMOS_VTL L=5e-08 W=9e-08 AD=5.175e-14 AS=5.175e-14 PD=1.33e-06 PS=1.33e-06 $X=59565 $Y=8195 $D=1
M194 186 B<12> gnd! gnd! NMOS_VTL L=5e-08 W=9e-08 AD=5.175e-14 AS=5.175e-14 PD=1.33e-06 PS=1.33e-06 $X=59565 $Y=15595 $D=1
M195 187 B<14> gnd! gnd! NMOS_VTL L=5e-08 W=9e-08 AD=5.175e-14 AS=5.175e-14 PD=1.33e-06 PS=1.33e-06 $X=59565 $Y=22995 $D=1
M196 188 91 gnd! gnd! NMOS_VTL L=5e-08 W=9e-08 AD=5.175e-14 AS=5.175e-14 PD=1.33e-06 PS=1.33e-06 $X=63450 $Y=790 $D=1
M197 189 92 gnd! gnd! NMOS_VTL L=5e-08 W=9e-08 AD=5.175e-14 AS=5.175e-14 PD=1.33e-06 PS=1.33e-06 $X=63450 $Y=8190 $D=1
M198 190 93 gnd! gnd! NMOS_VTL L=5e-08 W=9e-08 AD=5.175e-14 AS=5.175e-14 PD=1.33e-06 PS=1.33e-06 $X=63450 $Y=15590 $D=1
M199 191 94 gnd! gnd! NMOS_VTL L=5e-08 W=9e-08 AD=5.175e-14 AS=5.175e-14 PD=1.33e-06 PS=1.33e-06 $X=63450 $Y=22990 $D=1
M200 Sout<9> 95 107 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.161e-13 AS=1.26e-13 PD=1.65e-06 PS=1.76e-06 $X=64000 $Y=6470 $D=1
M201 Sout<11> 96 108 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.161e-13 AS=1.26e-13 PD=1.65e-06 PS=1.76e-06 $X=64000 $Y=13870 $D=1
M202 Sout<13> 97 109 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.161e-13 AS=1.26e-13 PD=1.65e-06 PS=1.76e-06 $X=64000 $Y=21270 $D=1
M203 Sout<15> 98 110 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.161e-13 AS=1.26e-13 PD=1.65e-06 PS=1.76e-06 $X=64000 $Y=28670 $D=1
M204 332 192 Sout<9> gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=9.855e-14 AS=1.161e-13 PD=1.455e-06 PS=1.65e-06 $X=65390 $Y=6470 $D=1
M205 333 193 Sout<11> gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=9.855e-14 AS=1.161e-13 PD=1.455e-06 PS=1.65e-06 $X=65390 $Y=13870 $D=1
M206 334 194 Sout<13> gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=9.855e-14 AS=1.161e-13 PD=1.455e-06 PS=1.65e-06 $X=65390 $Y=21270 $D=1
M207 335 195 Sout<15> gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=9.855e-14 AS=1.161e-13 PD=1.455e-06 PS=1.65e-06 $X=65390 $Y=28670 $D=1
M208 gnd! 180 332 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.2285e-13 AS=9.855e-14 PD=1.725e-06 PS=1.455e-06 $X=66585 $Y=6470 $D=1
M209 gnd! 181 333 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.2285e-13 AS=9.855e-14 PD=1.725e-06 PS=1.455e-06 $X=66585 $Y=13870 $D=1
M210 gnd! 182 334 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.2285e-13 AS=9.855e-14 PD=1.725e-06 PS=1.455e-06 $X=66585 $Y=21270 $D=1
M211 gnd! 183 335 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.2285e-13 AS=9.855e-14 PD=1.725e-06 PS=1.455e-06 $X=66585 $Y=28670 $D=1
M212 gnd! 91 115 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.2285e-13 AS=4.05e-14 PD=1.725e-06 PS=8.1e-07 $X=66850 $Y=900 $D=1
M213 gnd! 92 116 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.2285e-13 AS=4.05e-14 PD=1.725e-06 PS=8.1e-07 $X=66850 $Y=8300 $D=1
M214 gnd! 93 117 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.2285e-13 AS=4.05e-14 PD=1.725e-06 PS=8.1e-07 $X=66850 $Y=15700 $D=1
M215 gnd! 94 118 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.2285e-13 AS=4.05e-14 PD=1.725e-06 PS=8.1e-07 $X=66850 $Y=23100 $D=1
M216 107 99 gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=4.05e-14 AS=1.2285e-13 PD=8.1e-07 PS=1.725e-06 $X=68050 $Y=6470 $D=1
M217 108 100 gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=4.05e-14 AS=1.2285e-13 PD=8.1e-07 PS=1.725e-06 $X=68050 $Y=13870 $D=1
M218 109 101 gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=4.05e-14 AS=1.2285e-13 PD=8.1e-07 PS=1.725e-06 $X=68050 $Y=21270 $D=1
M219 110 102 gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=4.05e-14 AS=1.2285e-13 PD=8.1e-07 PS=1.725e-06 $X=68050 $Y=28670 $D=1
M220 336 200 gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=9.855e-14 AS=1.2285e-13 PD=1.455e-06 PS=1.725e-06 $X=68315 $Y=900 $D=1
M221 337 201 gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=9.855e-14 AS=1.2285e-13 PD=1.455e-06 PS=1.725e-06 $X=68315 $Y=8300 $D=1
M222 338 202 gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=9.855e-14 AS=1.2285e-13 PD=1.455e-06 PS=1.725e-06 $X=68315 $Y=15700 $D=1
M223 339 203 gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=9.855e-14 AS=1.2285e-13 PD=1.455e-06 PS=1.725e-06 $X=68315 $Y=23100 $D=1
M224 Sout<8> 188 336 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.161e-13 AS=9.855e-14 PD=1.65e-06 PS=1.455e-06 $X=69510 $Y=900 $D=1
M225 Sout<10> 189 337 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.161e-13 AS=9.855e-14 PD=1.65e-06 PS=1.455e-06 $X=69510 $Y=8300 $D=1
M226 Sout<12> 190 338 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.161e-13 AS=9.855e-14 PD=1.65e-06 PS=1.455e-06 $X=69510 $Y=15700 $D=1
M227 Sout<14> 191 339 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.161e-13 AS=9.855e-14 PD=1.65e-06 PS=1.455e-06 $X=69510 $Y=23100 $D=1
M228 115 19 Sout<8> gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.26e-13 AS=1.161e-13 PD=1.76e-06 PS=1.65e-06 $X=70900 $Y=900 $D=1
M229 116 85 Sout<10> gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.26e-13 AS=1.161e-13 PD=1.76e-06 PS=1.65e-06 $X=70900 $Y=8300 $D=1
M230 117 84 Sout<12> gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.26e-13 AS=1.161e-13 PD=1.76e-06 PS=1.65e-06 $X=70900 $Y=15700 $D=1
M231 118 86 Sout<14> gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.26e-13 AS=1.161e-13 PD=1.76e-06 PS=1.65e-06 $X=70900 $Y=23100 $D=1
M232 gnd! 99 192 gnd! NMOS_VTL L=5e-08 W=9e-08 AD=5.175e-14 AS=5.175e-14 PD=1.33e-06 PS=1.33e-06 $X=71450 $Y=6760 $D=1
M233 gnd! 100 193 gnd! NMOS_VTL L=5e-08 W=9e-08 AD=5.175e-14 AS=5.175e-14 PD=1.33e-06 PS=1.33e-06 $X=71450 $Y=14160 $D=1
M234 gnd! 101 194 gnd! NMOS_VTL L=5e-08 W=9e-08 AD=5.175e-14 AS=5.175e-14 PD=1.33e-06 PS=1.33e-06 $X=71450 $Y=21560 $D=1
M235 gnd! 102 195 gnd! NMOS_VTL L=5e-08 W=9e-08 AD=5.175e-14 AS=5.175e-14 PD=1.33e-06 PS=1.33e-06 $X=71450 $Y=28960 $D=1
M236 gnd! B<9> 196 gnd! NMOS_VTL L=5e-08 W=9e-08 AD=5.175e-14 AS=5.175e-14 PD=1.33e-06 PS=1.33e-06 $X=75335 $Y=6755 $D=1
M237 gnd! B<11> 197 gnd! NMOS_VTL L=5e-08 W=9e-08 AD=5.175e-14 AS=5.175e-14 PD=1.33e-06 PS=1.33e-06 $X=75335 $Y=14155 $D=1
M238 gnd! B<13> 198 gnd! NMOS_VTL L=5e-08 W=9e-08 AD=5.175e-14 AS=5.175e-14 PD=1.33e-06 PS=1.33e-06 $X=75335 $Y=21555 $D=1
M239 gnd! B<15> 199 gnd! NMOS_VTL L=5e-08 W=9e-08 AD=5.175e-14 AS=5.175e-14 PD=1.33e-06 PS=1.33e-06 $X=75335 $Y=28955 $D=1
M240 200 19 gnd! gnd! NMOS_VTL L=5e-08 W=9e-08 AD=5.175e-14 AS=5.175e-14 PD=1.33e-06 PS=1.33e-06 $X=76065 $Y=795 $D=1
M241 201 85 gnd! gnd! NMOS_VTL L=5e-08 W=9e-08 AD=5.175e-14 AS=5.175e-14 PD=1.33e-06 PS=1.33e-06 $X=76065 $Y=8195 $D=1
M242 202 84 gnd! gnd! NMOS_VTL L=5e-08 W=9e-08 AD=5.175e-14 AS=5.175e-14 PD=1.33e-06 PS=1.33e-06 $X=76065 $Y=15595 $D=1
M243 203 86 gnd! gnd! NMOS_VTL L=5e-08 W=9e-08 AD=5.175e-14 AS=5.175e-14 PD=1.33e-06 PS=1.33e-06 $X=76065 $Y=22995 $D=1
M244 340 91 gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=8.82e-14 AS=7.155e-14 PD=1.34e-06 PS=1.155e-06 $X=79290 $Y=695 $D=1
M245 341 92 gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=8.82e-14 AS=7.155e-14 PD=1.34e-06 PS=1.155e-06 $X=79290 $Y=8095 $D=1
M246 342 93 gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=8.82e-14 AS=7.155e-14 PD=1.34e-06 PS=1.155e-06 $X=79290 $Y=15495 $D=1
M247 343 94 gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=8.82e-14 AS=7.155e-14 PD=1.34e-06 PS=1.155e-06 $X=79290 $Y=22895 $D=1
M248 204 19 340 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=8.595e-14 AS=8.82e-14 PD=1.315e-06 PS=1.34e-06 $X=80370 $Y=695 $D=1
M249 205 85 341 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=8.595e-14 AS=8.82e-14 PD=1.315e-06 PS=1.34e-06 $X=80370 $Y=8095 $D=1
M250 206 84 342 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=8.595e-14 AS=8.82e-14 PD=1.315e-06 PS=1.34e-06 $X=80370 $Y=15495 $D=1
M251 207 86 343 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=8.595e-14 AS=8.82e-14 PD=1.315e-06 PS=1.34e-06 $X=80370 $Y=22895 $D=1
M252 99 B<9> 123 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.161e-13 AS=1.26e-13 PD=1.65e-06 PS=1.76e-06 $X=80500 $Y=6470 $D=1
M253 100 B<11> 124 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.161e-13 AS=1.26e-13 PD=1.65e-06 PS=1.76e-06 $X=80500 $Y=13870 $D=1
M254 101 B<13> 125 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.161e-13 AS=1.26e-13 PD=1.65e-06 PS=1.76e-06 $X=80500 $Y=21270 $D=1
M255 102 B<15> 126 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.161e-13 AS=1.26e-13 PD=1.65e-06 PS=1.76e-06 $X=80500 $Y=28670 $D=1
M256 344 208 99 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=9.855e-14 AS=1.161e-13 PD=1.455e-06 PS=1.65e-06 $X=81890 $Y=6470 $D=1
M257 345 209 100 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=9.855e-14 AS=1.161e-13 PD=1.455e-06 PS=1.65e-06 $X=81890 $Y=13870 $D=1
M258 346 210 101 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=9.855e-14 AS=1.161e-13 PD=1.455e-06 PS=1.65e-06 $X=81890 $Y=21270 $D=1
M259 347 211 102 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=9.855e-14 AS=1.161e-13 PD=1.455e-06 PS=1.65e-06 $X=81890 $Y=28670 $D=1
M260 gnd! 196 344 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.2285e-13 AS=9.855e-14 PD=1.725e-06 PS=1.455e-06 $X=83085 $Y=6470 $D=1
M261 gnd! 197 345 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.2285e-13 AS=9.855e-14 PD=1.725e-06 PS=1.455e-06 $X=83085 $Y=13870 $D=1
M262 gnd! 198 346 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.2285e-13 AS=9.855e-14 PD=1.725e-06 PS=1.455e-06 $X=83085 $Y=21270 $D=1
M263 gnd! 199 347 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.2285e-13 AS=9.855e-14 PD=1.725e-06 PS=1.455e-06 $X=83085 $Y=28670 $D=1
M264 348 204 gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=8.82e-14 AS=7.155e-14 PD=1.34e-06 PS=1.155e-06 $X=83290 $Y=695 $D=1
M265 349 205 gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=8.82e-14 AS=7.155e-14 PD=1.34e-06 PS=1.155e-06 $X=83290 $Y=8095 $D=1
M266 350 206 gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=8.82e-14 AS=7.155e-14 PD=1.34e-06 PS=1.155e-06 $X=83290 $Y=15495 $D=1
M267 351 207 gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=8.82e-14 AS=7.155e-14 PD=1.34e-06 PS=1.155e-06 $X=83290 $Y=22895 $D=1
M268 95 127 348 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=8.595e-14 AS=8.82e-14 PD=1.315e-06 PS=1.34e-06 $X=84370 $Y=695 $D=1
M269 96 128 349 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=8.595e-14 AS=8.82e-14 PD=1.315e-06 PS=1.34e-06 $X=84370 $Y=8095 $D=1
M270 97 129 350 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=8.595e-14 AS=8.82e-14 PD=1.315e-06 PS=1.34e-06 $X=84370 $Y=15495 $D=1
M271 98 130 351 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=8.595e-14 AS=8.82e-14 PD=1.315e-06 PS=1.34e-06 $X=84370 $Y=22895 $D=1
M272 123 A<9> gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=4.05e-14 AS=1.2285e-13 PD=8.1e-07 PS=1.725e-06 $X=84550 $Y=6470 $D=1
M273 124 A<11> gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=4.05e-14 AS=1.2285e-13 PD=8.1e-07 PS=1.725e-06 $X=84550 $Y=13870 $D=1
M274 125 A<13> gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=4.05e-14 AS=1.2285e-13 PD=8.1e-07 PS=1.725e-06 $X=84550 $Y=21270 $D=1
M275 126 A<15> gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=4.05e-14 AS=1.2285e-13 PD=8.1e-07 PS=1.725e-06 $X=84550 $Y=28670 $D=1
M276 352 A<8> gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=8.82e-14 AS=7.155e-14 PD=1.34e-06 PS=1.155e-06 $X=87290 $Y=695 $D=1
M277 353 A<10> gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=8.82e-14 AS=7.155e-14 PD=1.34e-06 PS=1.155e-06 $X=87290 $Y=8095 $D=1
M278 354 A<12> gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=8.82e-14 AS=7.155e-14 PD=1.34e-06 PS=1.155e-06 $X=87290 $Y=15495 $D=1
M279 355 A<14> gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=8.82e-14 AS=7.155e-14 PD=1.34e-06 PS=1.155e-06 $X=87290 $Y=22895 $D=1
M280 gnd! A<9> 208 gnd! NMOS_VTL L=5e-08 W=9e-08 AD=5.175e-14 AS=5.175e-14 PD=1.33e-06 PS=1.33e-06 $X=87950 $Y=6760 $D=1
M281 gnd! A<11> 209 gnd! NMOS_VTL L=5e-08 W=9e-08 AD=5.175e-14 AS=5.175e-14 PD=1.33e-06 PS=1.33e-06 $X=87950 $Y=14160 $D=1
M282 gnd! A<13> 210 gnd! NMOS_VTL L=5e-08 W=9e-08 AD=5.175e-14 AS=5.175e-14 PD=1.33e-06 PS=1.33e-06 $X=87950 $Y=21560 $D=1
M283 gnd! A<15> 211 gnd! NMOS_VTL L=5e-08 W=9e-08 AD=5.175e-14 AS=5.175e-14 PD=1.33e-06 PS=1.33e-06 $X=87950 $Y=28960 $D=1
M284 127 B<8> 352 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=8.595e-14 AS=8.82e-14 PD=1.315e-06 PS=1.34e-06 $X=88370 $Y=695 $D=1
M285 128 B<10> 353 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=8.595e-14 AS=8.82e-14 PD=1.315e-06 PS=1.34e-06 $X=88370 $Y=8095 $D=1
M286 129 B<12> 354 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=8.595e-14 AS=8.82e-14 PD=1.315e-06 PS=1.34e-06 $X=88370 $Y=15495 $D=1
M287 130 B<14> 355 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=8.595e-14 AS=8.82e-14 PD=1.315e-06 PS=1.34e-06 $X=88370 $Y=22895 $D=1
M288 6 B<1> vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.65375e-13 AS=1.51031e-13 PD=1.655e-06 PS=1.57e-06 $X=1530 $Y=4490 $D=0
M289 7 B<3> vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.65375e-13 AS=1.51031e-13 PD=1.655e-06 PS=1.57e-06 $X=1530 $Y=11890 $D=0
M290 8 B<5> vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.65375e-13 AS=1.51031e-13 PD=1.655e-06 PS=1.57e-06 $X=1530 $Y=19290 $D=0
M291 9 B<7> vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.65375e-13 AS=1.51031e-13 PD=1.655e-06 PS=1.57e-06 $X=1530 $Y=26690 $D=0
M292 131 A<0> vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.94062e-13 AS=1.94062e-13 PD=1.825e-06 PS=1.825e-06 $X=1950 $Y=2630 $D=0
M293 132 A<2> vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.94062e-13 AS=1.94062e-13 PD=1.825e-06 PS=1.825e-06 $X=1950 $Y=10030 $D=0
M294 133 A<4> vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.94062e-13 AS=1.94062e-13 PD=1.825e-06 PS=1.825e-06 $X=1950 $Y=17430 $D=0
M295 134 A<6> vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.94062e-13 AS=1.94062e-13 PD=1.825e-06 PS=1.825e-06 $X=1950 $Y=24830 $D=0
M296 vdd! A<1> 6 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.34156e-13 AS=1.65375e-13 PD=1.47e-06 PS=1.655e-06 $X=2610 $Y=4490 $D=0
M297 vdd! A<3> 7 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.34156e-13 AS=1.65375e-13 PD=1.47e-06 PS=1.655e-06 $X=2610 $Y=11890 $D=0
M298 vdd! A<5> 8 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.34156e-13 AS=1.65375e-13 PD=1.47e-06 PS=1.655e-06 $X=2610 $Y=19290 $D=0
M299 vdd! A<7> 9 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.34156e-13 AS=1.65375e-13 PD=1.47e-06 PS=1.655e-06 $X=2610 $Y=26690 $D=0
M300 212 A<0> vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.30344e-13 AS=7.59375e-14 PD=2.04e-06 PS=1.125e-06 $X=5350 $Y=2565 $D=0
M301 213 A<2> vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.30344e-13 AS=7.59375e-14 PD=2.04e-06 PS=1.125e-06 $X=5350 $Y=9965 $D=0
M302 214 A<4> vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.30344e-13 AS=7.59375e-14 PD=2.04e-06 PS=1.125e-06 $X=5350 $Y=17365 $D=0
M303 215 A<6> vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.30344e-13 AS=7.59375e-14 PD=2.04e-06 PS=1.125e-06 $X=5350 $Y=24765 $D=0
M304 20 6 vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.65375e-13 AS=1.51031e-13 PD=1.655e-06 PS=1.57e-06 $X=5530 $Y=4490 $D=0
M305 18 7 vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.65375e-13 AS=1.51031e-13 PD=1.655e-06 PS=1.57e-06 $X=5530 $Y=11890 $D=0
M306 21 8 vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.65375e-13 AS=1.51031e-13 PD=1.655e-06 PS=1.57e-06 $X=5530 $Y=19290 $D=0
M307 19 9 vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.65375e-13 AS=1.51031e-13 PD=1.655e-06 PS=1.57e-06 $X=5530 $Y=26690 $D=0
M308 vdd! 135 20 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.34156e-13 AS=1.65375e-13 PD=1.47e-06 PS=1.655e-06 $X=6610 $Y=4490 $D=0
M309 vdd! 136 18 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.34156e-13 AS=1.65375e-13 PD=1.47e-06 PS=1.655e-06 $X=6610 $Y=11890 $D=0
M310 vdd! 137 21 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.34156e-13 AS=1.65375e-13 PD=1.47e-06 PS=1.655e-06 $X=6610 $Y=19290 $D=0
M311 vdd! 138 19 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.34156e-13 AS=1.65375e-13 PD=1.47e-06 PS=1.655e-06 $X=6610 $Y=26690 $D=0
M312 26 143 212 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.84781e-13 AS=2.30344e-13 PD=1.77e-06 PS=2.04e-06 $X=6815 $Y=2565 $D=0
M313 27 144 213 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.84781e-13 AS=2.30344e-13 PD=1.77e-06 PS=2.04e-06 $X=6815 $Y=9965 $D=0
M314 28 145 214 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.84781e-13 AS=2.30344e-13 PD=1.77e-06 PS=2.04e-06 $X=6815 $Y=17365 $D=0
M315 29 146 215 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.84781e-13 AS=2.30344e-13 PD=1.77e-06 PS=2.04e-06 $X=6815 $Y=24765 $D=0
M316 216 131 26 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.17687e-13 AS=1.84781e-13 PD=1.965e-06 PS=1.77e-06 $X=8010 $Y=2565 $D=0
M317 217 132 27 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.17687e-13 AS=1.84781e-13 PD=1.965e-06 PS=1.77e-06 $X=8010 $Y=9965 $D=0
M318 218 133 28 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.17687e-13 AS=1.84781e-13 PD=1.965e-06 PS=1.77e-06 $X=8010 $Y=17365 $D=0
M319 219 134 29 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.17687e-13 AS=1.84781e-13 PD=1.965e-06 PS=1.77e-06 $X=8010 $Y=24765 $D=0
M320 vdd! B<0> 216 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.3625e-13 AS=2.17687e-13 PD=2.075e-06 PS=1.965e-06 $X=9400 $Y=2565 $D=0
M321 vdd! B<2> 217 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.3625e-13 AS=2.17687e-13 PD=2.075e-06 PS=1.965e-06 $X=9400 $Y=9965 $D=0
M322 vdd! B<4> 218 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.3625e-13 AS=2.17687e-13 PD=2.075e-06 PS=1.965e-06 $X=9400 $Y=17365 $D=0
M323 vdd! B<6> 219 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.3625e-13 AS=2.17687e-13 PD=2.075e-06 PS=1.965e-06 $X=9400 $Y=24765 $D=0
M324 135 30 vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.65375e-13 AS=1.51031e-13 PD=1.655e-06 PS=1.57e-06 $X=9530 $Y=4490 $D=0
M325 136 31 vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.65375e-13 AS=1.51031e-13 PD=1.655e-06 PS=1.57e-06 $X=9530 $Y=11890 $D=0
M326 137 32 vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.65375e-13 AS=1.51031e-13 PD=1.655e-06 PS=1.57e-06 $X=9530 $Y=19290 $D=0
M327 138 33 vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.65375e-13 AS=1.51031e-13 PD=1.655e-06 PS=1.57e-06 $X=9530 $Y=26690 $D=0
M328 vdd! 34 135 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.34156e-13 AS=1.65375e-13 PD=1.47e-06 PS=1.655e-06 $X=10610 $Y=4490 $D=0
M329 vdd! 35 136 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.34156e-13 AS=1.65375e-13 PD=1.47e-06 PS=1.655e-06 $X=10610 $Y=11890 $D=0
M330 vdd! 36 137 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.34156e-13 AS=1.65375e-13 PD=1.47e-06 PS=1.655e-06 $X=10610 $Y=19290 $D=0
M331 vdd! 37 138 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.34156e-13 AS=1.65375e-13 PD=1.47e-06 PS=1.655e-06 $X=10610 $Y=26690 $D=0
M332 vdd! 30 139 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.94062e-13 AS=1.94062e-13 PD=1.825e-06 PS=1.825e-06 $X=13835 $Y=4420 $D=0
M333 vdd! 31 140 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.94062e-13 AS=1.94062e-13 PD=1.825e-06 PS=1.825e-06 $X=13835 $Y=11820 $D=0
M334 vdd! 32 141 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.94062e-13 AS=1.94062e-13 PD=1.825e-06 PS=1.825e-06 $X=13835 $Y=19220 $D=0
M335 vdd! 33 142 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.94062e-13 AS=1.94062e-13 PD=1.825e-06 PS=1.825e-06 $X=13835 $Y=26620 $D=0
M336 143 B<0> vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.94062e-13 AS=1.94062e-13 PD=1.825e-06 PS=1.825e-06 $X=14565 $Y=2635 $D=0
M337 144 B<2> vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.94062e-13 AS=1.94062e-13 PD=1.825e-06 PS=1.825e-06 $X=14565 $Y=10035 $D=0
M338 145 B<4> vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.94062e-13 AS=1.94062e-13 PD=1.825e-06 PS=1.825e-06 $X=14565 $Y=17435 $D=0
M339 146 B<6> vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.94062e-13 AS=1.94062e-13 PD=1.825e-06 PS=1.825e-06 $X=14565 $Y=24835 $D=0
M340 147 26 vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.94062e-13 AS=1.94062e-13 PD=1.825e-06 PS=1.825e-06 $X=18450 $Y=2630 $D=0
M341 148 27 vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.94062e-13 AS=1.94062e-13 PD=1.825e-06 PS=1.825e-06 $X=18450 $Y=10030 $D=0
M342 149 28 vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.94062e-13 AS=1.94062e-13 PD=1.825e-06 PS=1.825e-06 $X=18450 $Y=17430 $D=0
M343 150 29 vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.94062e-13 AS=1.94062e-13 PD=1.825e-06 PS=1.825e-06 $X=18450 $Y=24830 $D=0
M344 220 30 vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.17687e-13 AS=2.3625e-13 PD=1.965e-06 PS=2.075e-06 $X=19000 $Y=4490 $D=0
M345 221 31 vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.17687e-13 AS=2.3625e-13 PD=1.965e-06 PS=2.075e-06 $X=19000 $Y=11890 $D=0
M346 222 32 vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.17687e-13 AS=2.3625e-13 PD=1.965e-06 PS=2.075e-06 $X=19000 $Y=19290 $D=0
M347 223 33 vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.17687e-13 AS=2.3625e-13 PD=1.965e-06 PS=2.075e-06 $X=19000 $Y=26690 $D=0
M348 Sout<1> 151 220 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.84781e-13 AS=2.17687e-13 PD=1.77e-06 PS=1.965e-06 $X=20390 $Y=4490 $D=0
M349 Sout<3> 152 221 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.84781e-13 AS=2.17687e-13 PD=1.77e-06 PS=1.965e-06 $X=20390 $Y=11890 $D=0
M350 Sout<5> 153 222 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.84781e-13 AS=2.17687e-13 PD=1.77e-06 PS=1.965e-06 $X=20390 $Y=19290 $D=0
M351 Sout<7> 154 223 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.84781e-13 AS=2.17687e-13 PD=1.77e-06 PS=1.965e-06 $X=20390 $Y=26690 $D=0
M352 224 139 Sout<1> vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.30344e-13 AS=1.84781e-13 PD=2.04e-06 PS=1.77e-06 $X=21585 $Y=4490 $D=0
M353 225 140 Sout<3> vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.30344e-13 AS=1.84781e-13 PD=2.04e-06 PS=1.77e-06 $X=21585 $Y=11890 $D=0
M354 226 141 Sout<5> vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.30344e-13 AS=1.84781e-13 PD=2.04e-06 PS=1.77e-06 $X=21585 $Y=19290 $D=0
M355 227 142 Sout<7> vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.30344e-13 AS=1.84781e-13 PD=2.04e-06 PS=1.77e-06 $X=21585 $Y=26690 $D=0
M356 228 26 vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.30344e-13 AS=7.59375e-14 PD=2.04e-06 PS=1.125e-06 $X=21850 $Y=2565 $D=0
M357 229 27 vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.30344e-13 AS=7.59375e-14 PD=2.04e-06 PS=1.125e-06 $X=21850 $Y=9965 $D=0
M358 230 28 vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.30344e-13 AS=7.59375e-14 PD=2.04e-06 PS=1.125e-06 $X=21850 $Y=17365 $D=0
M359 231 29 vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.30344e-13 AS=7.59375e-14 PD=2.04e-06 PS=1.125e-06 $X=21850 $Y=24765 $D=0
M360 vdd! 34 224 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=7.59375e-14 AS=2.30344e-13 PD=1.125e-06 PS=2.04e-06 $X=23050 $Y=4490 $D=0
M361 vdd! 35 225 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=7.59375e-14 AS=2.30344e-13 PD=1.125e-06 PS=2.04e-06 $X=23050 $Y=11890 $D=0
M362 vdd! 36 226 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=7.59375e-14 AS=2.30344e-13 PD=1.125e-06 PS=2.04e-06 $X=23050 $Y=19290 $D=0
M363 vdd! 37 227 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=7.59375e-14 AS=2.30344e-13 PD=1.125e-06 PS=2.04e-06 $X=23050 $Y=26690 $D=0
M364 Sout<0> 159 228 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.84781e-13 AS=2.30344e-13 PD=1.77e-06 PS=2.04e-06 $X=23315 $Y=2565 $D=0
M365 Sout<2> 160 229 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.84781e-13 AS=2.30344e-13 PD=1.77e-06 PS=2.04e-06 $X=23315 $Y=9965 $D=0
M366 Sout<4> 161 230 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.84781e-13 AS=2.30344e-13 PD=1.77e-06 PS=2.04e-06 $X=23315 $Y=17365 $D=0
M367 Sout<6> 162 231 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.84781e-13 AS=2.30344e-13 PD=1.77e-06 PS=2.04e-06 $X=23315 $Y=24765 $D=0
M368 232 147 Sout<0> vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.17687e-13 AS=1.84781e-13 PD=1.965e-06 PS=1.77e-06 $X=24510 $Y=2565 $D=0
M369 233 148 Sout<2> vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.17687e-13 AS=1.84781e-13 PD=1.965e-06 PS=1.77e-06 $X=24510 $Y=9965 $D=0
M370 234 149 Sout<4> vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.17687e-13 AS=1.84781e-13 PD=1.965e-06 PS=1.77e-06 $X=24510 $Y=17365 $D=0
M371 235 150 Sout<6> vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.17687e-13 AS=1.84781e-13 PD=1.965e-06 PS=1.77e-06 $X=24510 $Y=24765 $D=0
M372 vdd! Cin 232 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.3625e-13 AS=2.17687e-13 PD=2.075e-06 PS=1.965e-06 $X=25900 $Y=2565 $D=0
M373 vdd! 20 233 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.3625e-13 AS=2.17687e-13 PD=2.075e-06 PS=1.965e-06 $X=25900 $Y=9965 $D=0
M374 vdd! 18 234 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.3625e-13 AS=2.17687e-13 PD=2.075e-06 PS=1.965e-06 $X=25900 $Y=17365 $D=0
M375 vdd! 21 235 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.3625e-13 AS=2.17687e-13 PD=2.075e-06 PS=1.965e-06 $X=25900 $Y=24765 $D=0
M376 vdd! 34 151 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.94062e-13 AS=1.94062e-13 PD=1.825e-06 PS=1.825e-06 $X=26450 $Y=4425 $D=0
M377 vdd! 35 152 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.94062e-13 AS=1.94062e-13 PD=1.825e-06 PS=1.825e-06 $X=26450 $Y=11825 $D=0
M378 vdd! 36 153 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.94062e-13 AS=1.94062e-13 PD=1.825e-06 PS=1.825e-06 $X=26450 $Y=19225 $D=0
M379 vdd! 37 154 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.94062e-13 AS=1.94062e-13 PD=1.825e-06 PS=1.825e-06 $X=26450 $Y=26625 $D=0
M380 vdd! B<1> 155 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.94062e-13 AS=1.94062e-13 PD=1.825e-06 PS=1.825e-06 $X=30335 $Y=4420 $D=0
M381 vdd! B<3> 156 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.94062e-13 AS=1.94062e-13 PD=1.825e-06 PS=1.825e-06 $X=30335 $Y=11820 $D=0
M382 vdd! B<5> 157 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.94062e-13 AS=1.94062e-13 PD=1.825e-06 PS=1.825e-06 $X=30335 $Y=19220 $D=0
M383 vdd! B<7> 158 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.94062e-13 AS=1.94062e-13 PD=1.825e-06 PS=1.825e-06 $X=30335 $Y=26620 $D=0
M384 159 Cin vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.94062e-13 AS=1.94062e-13 PD=1.825e-06 PS=1.825e-06 $X=31065 $Y=2635 $D=0
M385 160 20 vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.94062e-13 AS=1.94062e-13 PD=1.825e-06 PS=1.825e-06 $X=31065 $Y=10035 $D=0
M386 161 18 vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.94062e-13 AS=1.94062e-13 PD=1.825e-06 PS=1.825e-06 $X=31065 $Y=17435 $D=0
M387 162 21 vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.94062e-13 AS=1.94062e-13 PD=1.825e-06 PS=1.825e-06 $X=31065 $Y=24835 $D=0
M388 163 26 vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.65375e-13 AS=1.34156e-13 PD=1.655e-06 PS=1.47e-06 $X=34290 $Y=2565 $D=0
M389 164 27 vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.65375e-13 AS=1.34156e-13 PD=1.655e-06 PS=1.47e-06 $X=34290 $Y=9965 $D=0
M390 165 28 vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.65375e-13 AS=1.34156e-13 PD=1.655e-06 PS=1.47e-06 $X=34290 $Y=17365 $D=0
M391 166 29 vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.65375e-13 AS=1.34156e-13 PD=1.655e-06 PS=1.47e-06 $X=34290 $Y=24765 $D=0
M392 vdd! Cin 163 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.51031e-13 AS=1.65375e-13 PD=1.57e-06 PS=1.655e-06 $X=35370 $Y=2565 $D=0
M393 vdd! 20 164 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.51031e-13 AS=1.65375e-13 PD=1.57e-06 PS=1.655e-06 $X=35370 $Y=9965 $D=0
M394 vdd! 18 165 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.51031e-13 AS=1.65375e-13 PD=1.57e-06 PS=1.655e-06 $X=35370 $Y=17365 $D=0
M395 vdd! 21 166 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.51031e-13 AS=1.65375e-13 PD=1.57e-06 PS=1.655e-06 $X=35370 $Y=24765 $D=0
M396 236 B<1> vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.17687e-13 AS=2.3625e-13 PD=1.965e-06 PS=2.075e-06 $X=35500 $Y=4490 $D=0
M397 237 B<3> vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.17687e-13 AS=2.3625e-13 PD=1.965e-06 PS=2.075e-06 $X=35500 $Y=11890 $D=0
M398 238 B<5> vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.17687e-13 AS=2.3625e-13 PD=1.965e-06 PS=2.075e-06 $X=35500 $Y=19290 $D=0
M399 239 B<7> vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.17687e-13 AS=2.3625e-13 PD=1.965e-06 PS=2.075e-06 $X=35500 $Y=26690 $D=0
M400 34 167 236 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.84781e-13 AS=2.17687e-13 PD=1.77e-06 PS=1.965e-06 $X=36890 $Y=4490 $D=0
M401 35 168 237 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.84781e-13 AS=2.17687e-13 PD=1.77e-06 PS=1.965e-06 $X=36890 $Y=11890 $D=0
M402 36 169 238 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.84781e-13 AS=2.17687e-13 PD=1.77e-06 PS=1.965e-06 $X=36890 $Y=19290 $D=0
M403 37 170 239 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.84781e-13 AS=2.17687e-13 PD=1.77e-06 PS=1.965e-06 $X=36890 $Y=26690 $D=0
M404 240 155 34 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.30344e-13 AS=1.84781e-13 PD=2.04e-06 PS=1.77e-06 $X=38085 $Y=4490 $D=0
M405 241 156 35 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.30344e-13 AS=1.84781e-13 PD=2.04e-06 PS=1.77e-06 $X=38085 $Y=11890 $D=0
M406 242 157 36 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.30344e-13 AS=1.84781e-13 PD=2.04e-06 PS=1.77e-06 $X=38085 $Y=19290 $D=0
M407 243 158 37 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.30344e-13 AS=1.84781e-13 PD=2.04e-06 PS=1.77e-06 $X=38085 $Y=26690 $D=0
M408 30 163 vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.65375e-13 AS=1.34156e-13 PD=1.655e-06 PS=1.47e-06 $X=38290 $Y=2565 $D=0
M409 31 164 vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.65375e-13 AS=1.34156e-13 PD=1.655e-06 PS=1.47e-06 $X=38290 $Y=9965 $D=0
M410 32 165 vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.65375e-13 AS=1.34156e-13 PD=1.655e-06 PS=1.47e-06 $X=38290 $Y=17365 $D=0
M411 33 166 vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.65375e-13 AS=1.34156e-13 PD=1.655e-06 PS=1.47e-06 $X=38290 $Y=24765 $D=0
M412 vdd! 63 30 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.51031e-13 AS=1.65375e-13 PD=1.57e-06 PS=1.655e-06 $X=39370 $Y=2565 $D=0
M413 vdd! 64 31 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.51031e-13 AS=1.65375e-13 PD=1.57e-06 PS=1.655e-06 $X=39370 $Y=9965 $D=0
M414 vdd! 65 32 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.51031e-13 AS=1.65375e-13 PD=1.57e-06 PS=1.655e-06 $X=39370 $Y=17365 $D=0
M415 vdd! 66 33 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.51031e-13 AS=1.65375e-13 PD=1.57e-06 PS=1.655e-06 $X=39370 $Y=24765 $D=0
M416 vdd! A<1> 240 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=7.59375e-14 AS=2.30344e-13 PD=1.125e-06 PS=2.04e-06 $X=39550 $Y=4490 $D=0
M417 vdd! A<3> 241 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=7.59375e-14 AS=2.30344e-13 PD=1.125e-06 PS=2.04e-06 $X=39550 $Y=11890 $D=0
M418 vdd! A<5> 242 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=7.59375e-14 AS=2.30344e-13 PD=1.125e-06 PS=2.04e-06 $X=39550 $Y=19290 $D=0
M419 vdd! A<7> 243 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=7.59375e-14 AS=2.30344e-13 PD=1.125e-06 PS=2.04e-06 $X=39550 $Y=26690 $D=0
M420 63 A<0> vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.65375e-13 AS=1.34156e-13 PD=1.655e-06 PS=1.47e-06 $X=42290 $Y=2565 $D=0
M421 64 A<2> vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.65375e-13 AS=1.34156e-13 PD=1.655e-06 PS=1.47e-06 $X=42290 $Y=9965 $D=0
M422 65 A<4> vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.65375e-13 AS=1.34156e-13 PD=1.655e-06 PS=1.47e-06 $X=42290 $Y=17365 $D=0
M423 66 A<6> vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.65375e-13 AS=1.34156e-13 PD=1.655e-06 PS=1.47e-06 $X=42290 $Y=24765 $D=0
M424 vdd! A<1> 167 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.94062e-13 AS=1.94062e-13 PD=1.825e-06 PS=1.825e-06 $X=42950 $Y=4425 $D=0
M425 vdd! A<3> 168 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.94062e-13 AS=1.94062e-13 PD=1.825e-06 PS=1.825e-06 $X=42950 $Y=11825 $D=0
M426 vdd! A<5> 169 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.94062e-13 AS=1.94062e-13 PD=1.825e-06 PS=1.825e-06 $X=42950 $Y=19225 $D=0
M427 vdd! A<7> 170 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.94062e-13 AS=1.94062e-13 PD=1.825e-06 PS=1.825e-06 $X=42950 $Y=26625 $D=0
M428 vdd! B<0> 63 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.51031e-13 AS=1.65375e-13 PD=1.57e-06 PS=1.655e-06 $X=43370 $Y=2565 $D=0
M429 vdd! B<2> 64 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.51031e-13 AS=1.65375e-13 PD=1.57e-06 PS=1.655e-06 $X=43370 $Y=9965 $D=0
M430 vdd! B<4> 65 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.51031e-13 AS=1.65375e-13 PD=1.57e-06 PS=1.655e-06 $X=43370 $Y=17365 $D=0
M431 vdd! B<6> 66 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.51031e-13 AS=1.65375e-13 PD=1.57e-06 PS=1.655e-06 $X=43370 $Y=24765 $D=0
M432 72 B<9> vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.65375e-13 AS=1.51031e-13 PD=1.655e-06 PS=1.57e-06 $X=46530 $Y=4490 $D=0
M433 73 B<11> vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.65375e-13 AS=1.51031e-13 PD=1.655e-06 PS=1.57e-06 $X=46530 $Y=11890 $D=0
M434 74 B<13> vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.65375e-13 AS=1.51031e-13 PD=1.655e-06 PS=1.57e-06 $X=46530 $Y=19290 $D=0
M435 75 B<15> vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.65375e-13 AS=1.51031e-13 PD=1.655e-06 PS=1.57e-06 $X=46530 $Y=26690 $D=0
M436 171 A<8> vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.94062e-13 AS=1.94062e-13 PD=1.825e-06 PS=1.825e-06 $X=46950 $Y=2630 $D=0
M437 172 A<10> vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.94062e-13 AS=1.94062e-13 PD=1.825e-06 PS=1.825e-06 $X=46950 $Y=10030 $D=0
M438 173 A<12> vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.94062e-13 AS=1.94062e-13 PD=1.825e-06 PS=1.825e-06 $X=46950 $Y=17430 $D=0
M439 174 A<14> vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.94062e-13 AS=1.94062e-13 PD=1.825e-06 PS=1.825e-06 $X=46950 $Y=24830 $D=0
M440 vdd! A<9> 72 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.34156e-13 AS=1.65375e-13 PD=1.47e-06 PS=1.655e-06 $X=47610 $Y=4490 $D=0
M441 vdd! A<11> 73 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.34156e-13 AS=1.65375e-13 PD=1.47e-06 PS=1.655e-06 $X=47610 $Y=11890 $D=0
M442 vdd! A<13> 74 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.34156e-13 AS=1.65375e-13 PD=1.47e-06 PS=1.655e-06 $X=47610 $Y=19290 $D=0
M443 vdd! A<15> 75 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.34156e-13 AS=1.65375e-13 PD=1.47e-06 PS=1.655e-06 $X=47610 $Y=26690 $D=0
M444 244 A<8> vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.30344e-13 AS=7.59375e-14 PD=2.04e-06 PS=1.125e-06 $X=50350 $Y=2565 $D=0
M445 245 A<10> vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.30344e-13 AS=7.59375e-14 PD=2.04e-06 PS=1.125e-06 $X=50350 $Y=9965 $D=0
M446 246 A<12> vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.30344e-13 AS=7.59375e-14 PD=2.04e-06 PS=1.125e-06 $X=50350 $Y=17365 $D=0
M447 247 A<14> vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.30344e-13 AS=7.59375e-14 PD=2.04e-06 PS=1.125e-06 $X=50350 $Y=24765 $D=0
M448 85 72 vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.65375e-13 AS=1.51031e-13 PD=1.655e-06 PS=1.57e-06 $X=50530 $Y=4490 $D=0
M449 84 73 vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.65375e-13 AS=1.51031e-13 PD=1.655e-06 PS=1.57e-06 $X=50530 $Y=11890 $D=0
M450 86 74 vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.65375e-13 AS=1.51031e-13 PD=1.655e-06 PS=1.57e-06 $X=50530 $Y=19290 $D=0
M451 Cout 75 vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.65375e-13 AS=1.51031e-13 PD=1.655e-06 PS=1.57e-06 $X=50530 $Y=26690 $D=0
M452 vdd! 176 85 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.34156e-13 AS=1.65375e-13 PD=1.47e-06 PS=1.655e-06 $X=51610 $Y=4490 $D=0
M453 vdd! 177 84 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.34156e-13 AS=1.65375e-13 PD=1.47e-06 PS=1.655e-06 $X=51610 $Y=11890 $D=0
M454 vdd! 178 86 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.34156e-13 AS=1.65375e-13 PD=1.47e-06 PS=1.655e-06 $X=51610 $Y=19290 $D=0
M455 vdd! 179 Cout vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.34156e-13 AS=1.65375e-13 PD=1.47e-06 PS=1.655e-06 $X=51610 $Y=26690 $D=0
M456 91 184 244 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.84781e-13 AS=2.30344e-13 PD=1.77e-06 PS=2.04e-06 $X=51815 $Y=2565 $D=0
M457 92 185 245 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.84781e-13 AS=2.30344e-13 PD=1.77e-06 PS=2.04e-06 $X=51815 $Y=9965 $D=0
M458 93 186 246 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.84781e-13 AS=2.30344e-13 PD=1.77e-06 PS=2.04e-06 $X=51815 $Y=17365 $D=0
M459 94 187 247 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.84781e-13 AS=2.30344e-13 PD=1.77e-06 PS=2.04e-06 $X=51815 $Y=24765 $D=0
M460 248 171 91 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.17687e-13 AS=1.84781e-13 PD=1.965e-06 PS=1.77e-06 $X=53010 $Y=2565 $D=0
M461 249 172 92 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.17687e-13 AS=1.84781e-13 PD=1.965e-06 PS=1.77e-06 $X=53010 $Y=9965 $D=0
M462 250 173 93 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.17687e-13 AS=1.84781e-13 PD=1.965e-06 PS=1.77e-06 $X=53010 $Y=17365 $D=0
M463 251 174 94 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.17687e-13 AS=1.84781e-13 PD=1.965e-06 PS=1.77e-06 $X=53010 $Y=24765 $D=0
M464 vdd! B<8> 248 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.3625e-13 AS=2.17687e-13 PD=2.075e-06 PS=1.965e-06 $X=54400 $Y=2565 $D=0
M465 vdd! B<10> 249 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.3625e-13 AS=2.17687e-13 PD=2.075e-06 PS=1.965e-06 $X=54400 $Y=9965 $D=0
M466 vdd! B<12> 250 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.3625e-13 AS=2.17687e-13 PD=2.075e-06 PS=1.965e-06 $X=54400 $Y=17365 $D=0
M467 vdd! B<14> 251 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.3625e-13 AS=2.17687e-13 PD=2.075e-06 PS=1.965e-06 $X=54400 $Y=24765 $D=0
M468 176 95 vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.65375e-13 AS=1.51031e-13 PD=1.655e-06 PS=1.57e-06 $X=54530 $Y=4490 $D=0
M469 177 96 vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.65375e-13 AS=1.51031e-13 PD=1.655e-06 PS=1.57e-06 $X=54530 $Y=11890 $D=0
M470 178 97 vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.65375e-13 AS=1.51031e-13 PD=1.655e-06 PS=1.57e-06 $X=54530 $Y=19290 $D=0
M471 179 98 vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.65375e-13 AS=1.51031e-13 PD=1.655e-06 PS=1.57e-06 $X=54530 $Y=26690 $D=0
M472 vdd! 99 176 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.34156e-13 AS=1.65375e-13 PD=1.47e-06 PS=1.655e-06 $X=55610 $Y=4490 $D=0
M473 vdd! 100 177 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.34156e-13 AS=1.65375e-13 PD=1.47e-06 PS=1.655e-06 $X=55610 $Y=11890 $D=0
M474 vdd! 101 178 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.34156e-13 AS=1.65375e-13 PD=1.47e-06 PS=1.655e-06 $X=55610 $Y=19290 $D=0
M475 vdd! 102 179 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.34156e-13 AS=1.65375e-13 PD=1.47e-06 PS=1.655e-06 $X=55610 $Y=26690 $D=0
M476 vdd! 95 180 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.94062e-13 AS=1.94062e-13 PD=1.825e-06 PS=1.825e-06 $X=58835 $Y=4420 $D=0
M477 vdd! 96 181 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.94062e-13 AS=1.94062e-13 PD=1.825e-06 PS=1.825e-06 $X=58835 $Y=11820 $D=0
M478 vdd! 97 182 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.94062e-13 AS=1.94062e-13 PD=1.825e-06 PS=1.825e-06 $X=58835 $Y=19220 $D=0
M479 vdd! 98 183 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.94062e-13 AS=1.94062e-13 PD=1.825e-06 PS=1.825e-06 $X=58835 $Y=26620 $D=0
M480 184 B<8> vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.94062e-13 AS=1.94062e-13 PD=1.825e-06 PS=1.825e-06 $X=59565 $Y=2635 $D=0
M481 185 B<10> vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.94062e-13 AS=1.94062e-13 PD=1.825e-06 PS=1.825e-06 $X=59565 $Y=10035 $D=0
M482 186 B<12> vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.94062e-13 AS=1.94062e-13 PD=1.825e-06 PS=1.825e-06 $X=59565 $Y=17435 $D=0
M483 187 B<14> vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.94062e-13 AS=1.94062e-13 PD=1.825e-06 PS=1.825e-06 $X=59565 $Y=24835 $D=0
M484 188 91 vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.94062e-13 AS=1.94062e-13 PD=1.825e-06 PS=1.825e-06 $X=63450 $Y=2630 $D=0
M485 189 92 vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.94062e-13 AS=1.94062e-13 PD=1.825e-06 PS=1.825e-06 $X=63450 $Y=10030 $D=0
M486 190 93 vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.94062e-13 AS=1.94062e-13 PD=1.825e-06 PS=1.825e-06 $X=63450 $Y=17430 $D=0
M487 191 94 vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.94062e-13 AS=1.94062e-13 PD=1.825e-06 PS=1.825e-06 $X=63450 $Y=24830 $D=0
M488 252 95 vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.17687e-13 AS=2.3625e-13 PD=1.965e-06 PS=2.075e-06 $X=64000 $Y=4490 $D=0
M489 253 96 vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.17687e-13 AS=2.3625e-13 PD=1.965e-06 PS=2.075e-06 $X=64000 $Y=11890 $D=0
M490 254 97 vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.17687e-13 AS=2.3625e-13 PD=1.965e-06 PS=2.075e-06 $X=64000 $Y=19290 $D=0
M491 255 98 vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.17687e-13 AS=2.3625e-13 PD=1.965e-06 PS=2.075e-06 $X=64000 $Y=26690 $D=0
M492 Sout<9> 192 252 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.84781e-13 AS=2.17687e-13 PD=1.77e-06 PS=1.965e-06 $X=65390 $Y=4490 $D=0
M493 Sout<11> 193 253 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.84781e-13 AS=2.17687e-13 PD=1.77e-06 PS=1.965e-06 $X=65390 $Y=11890 $D=0
M494 Sout<13> 194 254 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.84781e-13 AS=2.17687e-13 PD=1.77e-06 PS=1.965e-06 $X=65390 $Y=19290 $D=0
M495 Sout<15> 195 255 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.84781e-13 AS=2.17687e-13 PD=1.77e-06 PS=1.965e-06 $X=65390 $Y=26690 $D=0
M496 256 180 Sout<9> vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.30344e-13 AS=1.84781e-13 PD=2.04e-06 PS=1.77e-06 $X=66585 $Y=4490 $D=0
M497 257 181 Sout<11> vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.30344e-13 AS=1.84781e-13 PD=2.04e-06 PS=1.77e-06 $X=66585 $Y=11890 $D=0
M498 258 182 Sout<13> vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.30344e-13 AS=1.84781e-13 PD=2.04e-06 PS=1.77e-06 $X=66585 $Y=19290 $D=0
M499 259 183 Sout<15> vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.30344e-13 AS=1.84781e-13 PD=2.04e-06 PS=1.77e-06 $X=66585 $Y=26690 $D=0
M500 260 91 vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.30344e-13 AS=7.59375e-14 PD=2.04e-06 PS=1.125e-06 $X=66850 $Y=2565 $D=0
M501 261 92 vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.30344e-13 AS=7.59375e-14 PD=2.04e-06 PS=1.125e-06 $X=66850 $Y=9965 $D=0
M502 262 93 vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.30344e-13 AS=7.59375e-14 PD=2.04e-06 PS=1.125e-06 $X=66850 $Y=17365 $D=0
M503 263 94 vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.30344e-13 AS=7.59375e-14 PD=2.04e-06 PS=1.125e-06 $X=66850 $Y=24765 $D=0
M504 vdd! 99 256 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=7.59375e-14 AS=2.30344e-13 PD=1.125e-06 PS=2.04e-06 $X=68050 $Y=4490 $D=0
M505 vdd! 100 257 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=7.59375e-14 AS=2.30344e-13 PD=1.125e-06 PS=2.04e-06 $X=68050 $Y=11890 $D=0
M506 vdd! 101 258 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=7.59375e-14 AS=2.30344e-13 PD=1.125e-06 PS=2.04e-06 $X=68050 $Y=19290 $D=0
M507 vdd! 102 259 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=7.59375e-14 AS=2.30344e-13 PD=1.125e-06 PS=2.04e-06 $X=68050 $Y=26690 $D=0
M508 Sout<8> 200 260 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.84781e-13 AS=2.30344e-13 PD=1.77e-06 PS=2.04e-06 $X=68315 $Y=2565 $D=0
M509 Sout<10> 201 261 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.84781e-13 AS=2.30344e-13 PD=1.77e-06 PS=2.04e-06 $X=68315 $Y=9965 $D=0
M510 Sout<12> 202 262 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.84781e-13 AS=2.30344e-13 PD=1.77e-06 PS=2.04e-06 $X=68315 $Y=17365 $D=0
M511 Sout<14> 203 263 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.84781e-13 AS=2.30344e-13 PD=1.77e-06 PS=2.04e-06 $X=68315 $Y=24765 $D=0
M512 264 188 Sout<8> vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.17687e-13 AS=1.84781e-13 PD=1.965e-06 PS=1.77e-06 $X=69510 $Y=2565 $D=0
M513 265 189 Sout<10> vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.17687e-13 AS=1.84781e-13 PD=1.965e-06 PS=1.77e-06 $X=69510 $Y=9965 $D=0
M514 266 190 Sout<12> vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.17687e-13 AS=1.84781e-13 PD=1.965e-06 PS=1.77e-06 $X=69510 $Y=17365 $D=0
M515 267 191 Sout<14> vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.17687e-13 AS=1.84781e-13 PD=1.965e-06 PS=1.77e-06 $X=69510 $Y=24765 $D=0
M516 vdd! 19 264 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.3625e-13 AS=2.17687e-13 PD=2.075e-06 PS=1.965e-06 $X=70900 $Y=2565 $D=0
M517 vdd! 85 265 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.3625e-13 AS=2.17687e-13 PD=2.075e-06 PS=1.965e-06 $X=70900 $Y=9965 $D=0
M518 vdd! 84 266 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.3625e-13 AS=2.17687e-13 PD=2.075e-06 PS=1.965e-06 $X=70900 $Y=17365 $D=0
M519 vdd! 86 267 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.3625e-13 AS=2.17687e-13 PD=2.075e-06 PS=1.965e-06 $X=70900 $Y=24765 $D=0
M520 vdd! 99 192 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.94062e-13 AS=1.94062e-13 PD=1.825e-06 PS=1.825e-06 $X=71450 $Y=4425 $D=0
M521 vdd! 100 193 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.94062e-13 AS=1.94062e-13 PD=1.825e-06 PS=1.825e-06 $X=71450 $Y=11825 $D=0
M522 vdd! 101 194 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.94062e-13 AS=1.94062e-13 PD=1.825e-06 PS=1.825e-06 $X=71450 $Y=19225 $D=0
M523 vdd! 102 195 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.94062e-13 AS=1.94062e-13 PD=1.825e-06 PS=1.825e-06 $X=71450 $Y=26625 $D=0
M524 vdd! B<9> 196 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.94062e-13 AS=1.94062e-13 PD=1.825e-06 PS=1.825e-06 $X=75335 $Y=4420 $D=0
M525 vdd! B<11> 197 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.94062e-13 AS=1.94062e-13 PD=1.825e-06 PS=1.825e-06 $X=75335 $Y=11820 $D=0
M526 vdd! B<13> 198 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.94062e-13 AS=1.94062e-13 PD=1.825e-06 PS=1.825e-06 $X=75335 $Y=19220 $D=0
M527 vdd! B<15> 199 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.94062e-13 AS=1.94062e-13 PD=1.825e-06 PS=1.825e-06 $X=75335 $Y=26620 $D=0
M528 200 19 vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.94062e-13 AS=1.94062e-13 PD=1.825e-06 PS=1.825e-06 $X=76065 $Y=2635 $D=0
M529 201 85 vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.94062e-13 AS=1.94062e-13 PD=1.825e-06 PS=1.825e-06 $X=76065 $Y=10035 $D=0
M530 202 84 vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.94062e-13 AS=1.94062e-13 PD=1.825e-06 PS=1.825e-06 $X=76065 $Y=17435 $D=0
M531 203 86 vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.94062e-13 AS=1.94062e-13 PD=1.825e-06 PS=1.825e-06 $X=76065 $Y=24835 $D=0
M532 204 91 vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.65375e-13 AS=1.34156e-13 PD=1.655e-06 PS=1.47e-06 $X=79290 $Y=2565 $D=0
M533 205 92 vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.65375e-13 AS=1.34156e-13 PD=1.655e-06 PS=1.47e-06 $X=79290 $Y=9965 $D=0
M534 206 93 vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.65375e-13 AS=1.34156e-13 PD=1.655e-06 PS=1.47e-06 $X=79290 $Y=17365 $D=0
M535 207 94 vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.65375e-13 AS=1.34156e-13 PD=1.655e-06 PS=1.47e-06 $X=79290 $Y=24765 $D=0
M536 vdd! 19 204 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.51031e-13 AS=1.65375e-13 PD=1.57e-06 PS=1.655e-06 $X=80370 $Y=2565 $D=0
M537 vdd! 85 205 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.51031e-13 AS=1.65375e-13 PD=1.57e-06 PS=1.655e-06 $X=80370 $Y=9965 $D=0
M538 vdd! 84 206 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.51031e-13 AS=1.65375e-13 PD=1.57e-06 PS=1.655e-06 $X=80370 $Y=17365 $D=0
M539 vdd! 86 207 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.51031e-13 AS=1.65375e-13 PD=1.57e-06 PS=1.655e-06 $X=80370 $Y=24765 $D=0
M540 268 B<9> vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.17687e-13 AS=2.3625e-13 PD=1.965e-06 PS=2.075e-06 $X=80500 $Y=4490 $D=0
M541 269 B<11> vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.17687e-13 AS=2.3625e-13 PD=1.965e-06 PS=2.075e-06 $X=80500 $Y=11890 $D=0
M542 270 B<13> vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.17687e-13 AS=2.3625e-13 PD=1.965e-06 PS=2.075e-06 $X=80500 $Y=19290 $D=0
M543 271 B<15> vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.17687e-13 AS=2.3625e-13 PD=1.965e-06 PS=2.075e-06 $X=80500 $Y=26690 $D=0
M544 99 208 268 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.84781e-13 AS=2.17687e-13 PD=1.77e-06 PS=1.965e-06 $X=81890 $Y=4490 $D=0
M545 100 209 269 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.84781e-13 AS=2.17687e-13 PD=1.77e-06 PS=1.965e-06 $X=81890 $Y=11890 $D=0
M546 101 210 270 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.84781e-13 AS=2.17687e-13 PD=1.77e-06 PS=1.965e-06 $X=81890 $Y=19290 $D=0
M547 102 211 271 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.84781e-13 AS=2.17687e-13 PD=1.77e-06 PS=1.965e-06 $X=81890 $Y=26690 $D=0
M548 272 196 99 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.30344e-13 AS=1.84781e-13 PD=2.04e-06 PS=1.77e-06 $X=83085 $Y=4490 $D=0
M549 273 197 100 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.30344e-13 AS=1.84781e-13 PD=2.04e-06 PS=1.77e-06 $X=83085 $Y=11890 $D=0
M550 274 198 101 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.30344e-13 AS=1.84781e-13 PD=2.04e-06 PS=1.77e-06 $X=83085 $Y=19290 $D=0
M551 275 199 102 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.30344e-13 AS=1.84781e-13 PD=2.04e-06 PS=1.77e-06 $X=83085 $Y=26690 $D=0
M552 95 204 vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.65375e-13 AS=1.34156e-13 PD=1.655e-06 PS=1.47e-06 $X=83290 $Y=2565 $D=0
M553 96 205 vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.65375e-13 AS=1.34156e-13 PD=1.655e-06 PS=1.47e-06 $X=83290 $Y=9965 $D=0
M554 97 206 vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.65375e-13 AS=1.34156e-13 PD=1.655e-06 PS=1.47e-06 $X=83290 $Y=17365 $D=0
M555 98 207 vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.65375e-13 AS=1.34156e-13 PD=1.655e-06 PS=1.47e-06 $X=83290 $Y=24765 $D=0
M556 vdd! 127 95 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.51031e-13 AS=1.65375e-13 PD=1.57e-06 PS=1.655e-06 $X=84370 $Y=2565 $D=0
M557 vdd! 128 96 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.51031e-13 AS=1.65375e-13 PD=1.57e-06 PS=1.655e-06 $X=84370 $Y=9965 $D=0
M558 vdd! 129 97 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.51031e-13 AS=1.65375e-13 PD=1.57e-06 PS=1.655e-06 $X=84370 $Y=17365 $D=0
M559 vdd! 130 98 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.51031e-13 AS=1.65375e-13 PD=1.57e-06 PS=1.655e-06 $X=84370 $Y=24765 $D=0
M560 vdd! A<9> 272 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=7.59375e-14 AS=2.30344e-13 PD=1.125e-06 PS=2.04e-06 $X=84550 $Y=4490 $D=0
M561 vdd! A<11> 273 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=7.59375e-14 AS=2.30344e-13 PD=1.125e-06 PS=2.04e-06 $X=84550 $Y=11890 $D=0
M562 vdd! A<13> 274 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=7.59375e-14 AS=2.30344e-13 PD=1.125e-06 PS=2.04e-06 $X=84550 $Y=19290 $D=0
M563 vdd! A<15> 275 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=7.59375e-14 AS=2.30344e-13 PD=1.125e-06 PS=2.04e-06 $X=84550 $Y=26690 $D=0
M564 127 A<8> vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.65375e-13 AS=1.34156e-13 PD=1.655e-06 PS=1.47e-06 $X=87290 $Y=2565 $D=0
M565 128 A<10> vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.65375e-13 AS=1.34156e-13 PD=1.655e-06 PS=1.47e-06 $X=87290 $Y=9965 $D=0
M566 129 A<12> vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.65375e-13 AS=1.34156e-13 PD=1.655e-06 PS=1.47e-06 $X=87290 $Y=17365 $D=0
M567 130 A<14> vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.65375e-13 AS=1.34156e-13 PD=1.655e-06 PS=1.47e-06 $X=87290 $Y=24765 $D=0
M568 vdd! A<9> 208 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.94062e-13 AS=1.94062e-13 PD=1.825e-06 PS=1.825e-06 $X=87950 $Y=4425 $D=0
M569 vdd! A<11> 209 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.94062e-13 AS=1.94062e-13 PD=1.825e-06 PS=1.825e-06 $X=87950 $Y=11825 $D=0
M570 vdd! A<13> 210 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.94062e-13 AS=1.94062e-13 PD=1.825e-06 PS=1.825e-06 $X=87950 $Y=19225 $D=0
M571 vdd! A<15> 211 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.94062e-13 AS=1.94062e-13 PD=1.825e-06 PS=1.825e-06 $X=87950 $Y=26625 $D=0
M572 vdd! B<8> 127 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.51031e-13 AS=1.65375e-13 PD=1.57e-06 PS=1.655e-06 $X=88370 $Y=2565 $D=0
M573 vdd! B<10> 128 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.51031e-13 AS=1.65375e-13 PD=1.57e-06 PS=1.655e-06 $X=88370 $Y=9965 $D=0
M574 vdd! B<12> 129 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.51031e-13 AS=1.65375e-13 PD=1.57e-06 PS=1.655e-06 $X=88370 $Y=17365 $D=0
M575 vdd! B<14> 130 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.51031e-13 AS=1.65375e-13 PD=1.57e-06 PS=1.655e-06 $X=88370 $Y=24765 $D=0
.ENDS
***************************************

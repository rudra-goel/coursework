* SPICE NETLIST
***************************************

.SUBCKT 4_bit_ripple_carry_adder gnd! B<1> B<3> A<0> A<2> A<1> A<3> B<0> B<2> Sout<1> Sout<3> Sout<0> Sout<2> C_in vdd! C_out
** N=91 EP=16 IP=0 FDC=144
M0 72 B<1> 4 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=8.82e-14 AS=8.595e-14 PD=1.34e-06 PS=1.315e-06 $X=1530 $Y=6675 $D=1
M1 73 B<3> 5 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=8.82e-14 AS=8.595e-14 PD=1.34e-06 PS=1.315e-06 $X=1530 $Y=14075 $D=1
M2 35 A<0> gnd! gnd! NMOS_VTL L=5e-08 W=9e-08 AD=5.175e-14 AS=5.175e-14 PD=1.33e-06 PS=1.33e-06 $X=1950 $Y=790 $D=1
M3 36 A<2> gnd! gnd! NMOS_VTL L=5e-08 W=9e-08 AD=5.175e-14 AS=5.175e-14 PD=1.33e-06 PS=1.33e-06 $X=1950 $Y=8190 $D=1
M4 gnd! A<1> 72 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=7.155e-14 AS=8.82e-14 PD=1.155e-06 PS=1.34e-06 $X=2610 $Y=6675 $D=1
M5 gnd! A<3> 73 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=7.155e-14 AS=8.82e-14 PD=1.155e-06 PS=1.34e-06 $X=2610 $Y=14075 $D=1
M6 gnd! A<0> 11 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.2285e-13 AS=4.05e-14 PD=1.725e-06 PS=8.1e-07 $X=5350 $Y=900 $D=1
M7 gnd! A<2> 12 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.2285e-13 AS=4.05e-14 PD=1.725e-06 PS=8.1e-07 $X=5350 $Y=8300 $D=1
M8 74 4 10 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=8.82e-14 AS=8.595e-14 PD=1.34e-06 PS=1.315e-06 $X=5530 $Y=6675 $D=1
M9 75 5 C_out gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=8.82e-14 AS=8.595e-14 PD=1.34e-06 PS=1.315e-06 $X=5530 $Y=14075 $D=1
M10 gnd! 38 74 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=7.155e-14 AS=8.82e-14 PD=1.155e-06 PS=1.34e-06 $X=6610 $Y=6675 $D=1
M11 gnd! 39 75 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=7.155e-14 AS=8.82e-14 PD=1.155e-06 PS=1.34e-06 $X=6610 $Y=14075 $D=1
M12 76 42 gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=9.855e-14 AS=1.2285e-13 PD=1.455e-06 PS=1.725e-06 $X=6815 $Y=900 $D=1
M13 77 43 gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=9.855e-14 AS=1.2285e-13 PD=1.455e-06 PS=1.725e-06 $X=6815 $Y=8300 $D=1
M14 13 35 76 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.161e-13 AS=9.855e-14 PD=1.65e-06 PS=1.455e-06 $X=8010 $Y=900 $D=1
M15 14 36 77 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.161e-13 AS=9.855e-14 PD=1.65e-06 PS=1.455e-06 $X=8010 $Y=8300 $D=1
M16 11 B<0> 13 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.26e-13 AS=1.161e-13 PD=1.76e-06 PS=1.65e-06 $X=9400 $Y=900 $D=1
M17 12 B<2> 14 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.26e-13 AS=1.161e-13 PD=1.76e-06 PS=1.65e-06 $X=9400 $Y=8300 $D=1
M18 78 15 38 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=8.82e-14 AS=8.595e-14 PD=1.34e-06 PS=1.315e-06 $X=9530 $Y=6675 $D=1
M19 79 16 39 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=8.82e-14 AS=8.595e-14 PD=1.34e-06 PS=1.315e-06 $X=9530 $Y=14075 $D=1
M20 gnd! 17 78 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=7.155e-14 AS=8.82e-14 PD=1.155e-06 PS=1.34e-06 $X=10610 $Y=6675 $D=1
M21 gnd! 18 79 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=7.155e-14 AS=8.82e-14 PD=1.155e-06 PS=1.34e-06 $X=10610 $Y=14075 $D=1
M22 gnd! 15 40 gnd! NMOS_VTL L=5e-08 W=9e-08 AD=5.175e-14 AS=5.175e-14 PD=1.33e-06 PS=1.33e-06 $X=13835 $Y=6755 $D=1
M23 gnd! 16 41 gnd! NMOS_VTL L=5e-08 W=9e-08 AD=5.175e-14 AS=5.175e-14 PD=1.33e-06 PS=1.33e-06 $X=13835 $Y=14155 $D=1
M24 42 B<0> gnd! gnd! NMOS_VTL L=5e-08 W=9e-08 AD=5.175e-14 AS=5.175e-14 PD=1.33e-06 PS=1.33e-06 $X=14565 $Y=795 $D=1
M25 43 B<2> gnd! gnd! NMOS_VTL L=5e-08 W=9e-08 AD=5.175e-14 AS=5.175e-14 PD=1.33e-06 PS=1.33e-06 $X=14565 $Y=8195 $D=1
M26 44 13 gnd! gnd! NMOS_VTL L=5e-08 W=9e-08 AD=5.175e-14 AS=5.175e-14 PD=1.33e-06 PS=1.33e-06 $X=18450 $Y=790 $D=1
M27 45 14 gnd! gnd! NMOS_VTL L=5e-08 W=9e-08 AD=5.175e-14 AS=5.175e-14 PD=1.33e-06 PS=1.33e-06 $X=18450 $Y=8190 $D=1
M28 Sout<1> 15 21 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.161e-13 AS=1.26e-13 PD=1.65e-06 PS=1.76e-06 $X=19000 $Y=6470 $D=1
M29 Sout<3> 16 22 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.161e-13 AS=1.26e-13 PD=1.65e-06 PS=1.76e-06 $X=19000 $Y=13870 $D=1
M30 80 46 Sout<1> gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=9.855e-14 AS=1.161e-13 PD=1.455e-06 PS=1.65e-06 $X=20390 $Y=6470 $D=1
M31 81 47 Sout<3> gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=9.855e-14 AS=1.161e-13 PD=1.455e-06 PS=1.65e-06 $X=20390 $Y=13870 $D=1
M32 gnd! 40 80 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.2285e-13 AS=9.855e-14 PD=1.725e-06 PS=1.455e-06 $X=21585 $Y=6470 $D=1
M33 gnd! 41 81 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.2285e-13 AS=9.855e-14 PD=1.725e-06 PS=1.455e-06 $X=21585 $Y=13870 $D=1
M34 gnd! 13 25 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.2285e-13 AS=4.05e-14 PD=1.725e-06 PS=8.1e-07 $X=21850 $Y=900 $D=1
M35 gnd! 14 26 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.2285e-13 AS=4.05e-14 PD=1.725e-06 PS=8.1e-07 $X=21850 $Y=8300 $D=1
M36 21 17 gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=4.05e-14 AS=1.2285e-13 PD=8.1e-07 PS=1.725e-06 $X=23050 $Y=6470 $D=1
M37 22 18 gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=4.05e-14 AS=1.2285e-13 PD=8.1e-07 PS=1.725e-06 $X=23050 $Y=13870 $D=1
M38 82 50 gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=9.855e-14 AS=1.2285e-13 PD=1.455e-06 PS=1.725e-06 $X=23315 $Y=900 $D=1
M39 83 51 gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=9.855e-14 AS=1.2285e-13 PD=1.455e-06 PS=1.725e-06 $X=23315 $Y=8300 $D=1
M40 Sout<0> 44 82 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.161e-13 AS=9.855e-14 PD=1.65e-06 PS=1.455e-06 $X=24510 $Y=900 $D=1
M41 Sout<2> 45 83 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.161e-13 AS=9.855e-14 PD=1.65e-06 PS=1.455e-06 $X=24510 $Y=8300 $D=1
M42 25 C_in Sout<0> gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.26e-13 AS=1.161e-13 PD=1.76e-06 PS=1.65e-06 $X=25900 $Y=900 $D=1
M43 26 10 Sout<2> gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.26e-13 AS=1.161e-13 PD=1.76e-06 PS=1.65e-06 $X=25900 $Y=8300 $D=1
M44 gnd! 17 46 gnd! NMOS_VTL L=5e-08 W=9e-08 AD=5.175e-14 AS=5.175e-14 PD=1.33e-06 PS=1.33e-06 $X=26450 $Y=6760 $D=1
M45 gnd! 18 47 gnd! NMOS_VTL L=5e-08 W=9e-08 AD=5.175e-14 AS=5.175e-14 PD=1.33e-06 PS=1.33e-06 $X=26450 $Y=14160 $D=1
M46 gnd! B<1> 48 gnd! NMOS_VTL L=5e-08 W=9e-08 AD=5.175e-14 AS=5.175e-14 PD=1.33e-06 PS=1.33e-06 $X=30335 $Y=6755 $D=1
M47 gnd! B<3> 49 gnd! NMOS_VTL L=5e-08 W=9e-08 AD=5.175e-14 AS=5.175e-14 PD=1.33e-06 PS=1.33e-06 $X=30335 $Y=14155 $D=1
M48 50 C_in gnd! gnd! NMOS_VTL L=5e-08 W=9e-08 AD=5.175e-14 AS=5.175e-14 PD=1.33e-06 PS=1.33e-06 $X=31065 $Y=795 $D=1
M49 51 10 gnd! gnd! NMOS_VTL L=5e-08 W=9e-08 AD=5.175e-14 AS=5.175e-14 PD=1.33e-06 PS=1.33e-06 $X=31065 $Y=8195 $D=1
M50 84 13 gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=8.82e-14 AS=7.155e-14 PD=1.34e-06 PS=1.155e-06 $X=34290 $Y=695 $D=1
M51 85 14 gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=8.82e-14 AS=7.155e-14 PD=1.34e-06 PS=1.155e-06 $X=34290 $Y=8095 $D=1
M52 52 C_in 84 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=8.595e-14 AS=8.82e-14 PD=1.315e-06 PS=1.34e-06 $X=35370 $Y=695 $D=1
M53 53 10 85 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=8.595e-14 AS=8.82e-14 PD=1.315e-06 PS=1.34e-06 $X=35370 $Y=8095 $D=1
M54 17 B<1> 30 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.161e-13 AS=1.26e-13 PD=1.65e-06 PS=1.76e-06 $X=35500 $Y=6470 $D=1
M55 18 B<3> 31 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.161e-13 AS=1.26e-13 PD=1.65e-06 PS=1.76e-06 $X=35500 $Y=13870 $D=1
M56 86 54 17 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=9.855e-14 AS=1.161e-13 PD=1.455e-06 PS=1.65e-06 $X=36890 $Y=6470 $D=1
M57 87 55 18 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=9.855e-14 AS=1.161e-13 PD=1.455e-06 PS=1.65e-06 $X=36890 $Y=13870 $D=1
M58 gnd! 48 86 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.2285e-13 AS=9.855e-14 PD=1.725e-06 PS=1.455e-06 $X=38085 $Y=6470 $D=1
M59 gnd! 49 87 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.2285e-13 AS=9.855e-14 PD=1.725e-06 PS=1.455e-06 $X=38085 $Y=13870 $D=1
M60 88 52 gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=8.82e-14 AS=7.155e-14 PD=1.34e-06 PS=1.155e-06 $X=38290 $Y=695 $D=1
M61 89 53 gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=8.82e-14 AS=7.155e-14 PD=1.34e-06 PS=1.155e-06 $X=38290 $Y=8095 $D=1
M62 15 32 88 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=8.595e-14 AS=8.82e-14 PD=1.315e-06 PS=1.34e-06 $X=39370 $Y=695 $D=1
M63 16 33 89 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=8.595e-14 AS=8.82e-14 PD=1.315e-06 PS=1.34e-06 $X=39370 $Y=8095 $D=1
M64 30 A<1> gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=4.05e-14 AS=1.2285e-13 PD=8.1e-07 PS=1.725e-06 $X=39550 $Y=6470 $D=1
M65 31 A<3> gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=4.05e-14 AS=1.2285e-13 PD=8.1e-07 PS=1.725e-06 $X=39550 $Y=13870 $D=1
M66 90 A<0> gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=8.82e-14 AS=7.155e-14 PD=1.34e-06 PS=1.155e-06 $X=42290 $Y=695 $D=1
M67 91 A<2> gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=8.82e-14 AS=7.155e-14 PD=1.34e-06 PS=1.155e-06 $X=42290 $Y=8095 $D=1
M68 gnd! A<1> 54 gnd! NMOS_VTL L=5e-08 W=9e-08 AD=5.175e-14 AS=5.175e-14 PD=1.33e-06 PS=1.33e-06 $X=42950 $Y=6760 $D=1
M69 gnd! A<3> 55 gnd! NMOS_VTL L=5e-08 W=9e-08 AD=5.175e-14 AS=5.175e-14 PD=1.33e-06 PS=1.33e-06 $X=42950 $Y=14160 $D=1
M70 32 B<0> 90 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=8.595e-14 AS=8.82e-14 PD=1.315e-06 PS=1.34e-06 $X=43370 $Y=695 $D=1
M71 33 B<2> 91 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=8.595e-14 AS=8.82e-14 PD=1.315e-06 PS=1.34e-06 $X=43370 $Y=8095 $D=1
M72 4 B<1> vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.65375e-13 AS=1.51031e-13 PD=1.655e-06 PS=1.57e-06 $X=1530 $Y=4490 $D=0
M73 5 B<3> vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.65375e-13 AS=1.51031e-13 PD=1.655e-06 PS=1.57e-06 $X=1530 $Y=11890 $D=0
M74 35 A<0> vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.94062e-13 AS=1.94062e-13 PD=1.825e-06 PS=1.825e-06 $X=1950 $Y=2630 $D=0
M75 36 A<2> vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.94062e-13 AS=1.94062e-13 PD=1.825e-06 PS=1.825e-06 $X=1950 $Y=10030 $D=0
M76 vdd! A<1> 4 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.34156e-13 AS=1.65375e-13 PD=1.47e-06 PS=1.655e-06 $X=2610 $Y=4490 $D=0
M77 vdd! A<3> 5 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.34156e-13 AS=1.65375e-13 PD=1.47e-06 PS=1.655e-06 $X=2610 $Y=11890 $D=0
M78 56 A<0> vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.30344e-13 AS=7.59375e-14 PD=2.04e-06 PS=1.125e-06 $X=5350 $Y=2565 $D=0
M79 57 A<2> vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.30344e-13 AS=7.59375e-14 PD=2.04e-06 PS=1.125e-06 $X=5350 $Y=9965 $D=0
M80 10 4 vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.65375e-13 AS=1.51031e-13 PD=1.655e-06 PS=1.57e-06 $X=5530 $Y=4490 $D=0
M81 C_out 5 vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.65375e-13 AS=1.51031e-13 PD=1.655e-06 PS=1.57e-06 $X=5530 $Y=11890 $D=0
M82 vdd! 38 10 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.34156e-13 AS=1.65375e-13 PD=1.47e-06 PS=1.655e-06 $X=6610 $Y=4490 $D=0
M83 vdd! 39 C_out vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.34156e-13 AS=1.65375e-13 PD=1.47e-06 PS=1.655e-06 $X=6610 $Y=11890 $D=0
M84 13 42 56 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.84781e-13 AS=2.30344e-13 PD=1.77e-06 PS=2.04e-06 $X=6815 $Y=2565 $D=0
M85 14 43 57 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.84781e-13 AS=2.30344e-13 PD=1.77e-06 PS=2.04e-06 $X=6815 $Y=9965 $D=0
M86 58 35 13 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.17687e-13 AS=1.84781e-13 PD=1.965e-06 PS=1.77e-06 $X=8010 $Y=2565 $D=0
M87 59 36 14 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.17687e-13 AS=1.84781e-13 PD=1.965e-06 PS=1.77e-06 $X=8010 $Y=9965 $D=0
M88 vdd! B<0> 58 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.3625e-13 AS=2.17687e-13 PD=2.075e-06 PS=1.965e-06 $X=9400 $Y=2565 $D=0
M89 vdd! B<2> 59 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.3625e-13 AS=2.17687e-13 PD=2.075e-06 PS=1.965e-06 $X=9400 $Y=9965 $D=0
M90 38 15 vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.65375e-13 AS=1.51031e-13 PD=1.655e-06 PS=1.57e-06 $X=9530 $Y=4490 $D=0
M91 39 16 vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.65375e-13 AS=1.51031e-13 PD=1.655e-06 PS=1.57e-06 $X=9530 $Y=11890 $D=0
M92 vdd! 17 38 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.34156e-13 AS=1.65375e-13 PD=1.47e-06 PS=1.655e-06 $X=10610 $Y=4490 $D=0
M93 vdd! 18 39 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.34156e-13 AS=1.65375e-13 PD=1.47e-06 PS=1.655e-06 $X=10610 $Y=11890 $D=0
M94 vdd! 15 40 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.94062e-13 AS=1.94062e-13 PD=1.825e-06 PS=1.825e-06 $X=13835 $Y=4420 $D=0
M95 vdd! 16 41 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.94062e-13 AS=1.94062e-13 PD=1.825e-06 PS=1.825e-06 $X=13835 $Y=11820 $D=0
M96 42 B<0> vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.94062e-13 AS=1.94062e-13 PD=1.825e-06 PS=1.825e-06 $X=14565 $Y=2635 $D=0
M97 43 B<2> vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.94062e-13 AS=1.94062e-13 PD=1.825e-06 PS=1.825e-06 $X=14565 $Y=10035 $D=0
M98 44 13 vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.94062e-13 AS=1.94062e-13 PD=1.825e-06 PS=1.825e-06 $X=18450 $Y=2630 $D=0
M99 45 14 vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.94062e-13 AS=1.94062e-13 PD=1.825e-06 PS=1.825e-06 $X=18450 $Y=10030 $D=0
M100 60 15 vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.17687e-13 AS=2.3625e-13 PD=1.965e-06 PS=2.075e-06 $X=19000 $Y=4490 $D=0
M101 61 16 vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.17687e-13 AS=2.3625e-13 PD=1.965e-06 PS=2.075e-06 $X=19000 $Y=11890 $D=0
M102 Sout<1> 46 60 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.84781e-13 AS=2.17687e-13 PD=1.77e-06 PS=1.965e-06 $X=20390 $Y=4490 $D=0
M103 Sout<3> 47 61 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.84781e-13 AS=2.17687e-13 PD=1.77e-06 PS=1.965e-06 $X=20390 $Y=11890 $D=0
M104 62 40 Sout<1> vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.30344e-13 AS=1.84781e-13 PD=2.04e-06 PS=1.77e-06 $X=21585 $Y=4490 $D=0
M105 63 41 Sout<3> vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.30344e-13 AS=1.84781e-13 PD=2.04e-06 PS=1.77e-06 $X=21585 $Y=11890 $D=0
M106 64 13 vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.30344e-13 AS=7.59375e-14 PD=2.04e-06 PS=1.125e-06 $X=21850 $Y=2565 $D=0
M107 65 14 vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.30344e-13 AS=7.59375e-14 PD=2.04e-06 PS=1.125e-06 $X=21850 $Y=9965 $D=0
M108 vdd! 17 62 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=7.59375e-14 AS=2.30344e-13 PD=1.125e-06 PS=2.04e-06 $X=23050 $Y=4490 $D=0
M109 vdd! 18 63 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=7.59375e-14 AS=2.30344e-13 PD=1.125e-06 PS=2.04e-06 $X=23050 $Y=11890 $D=0
M110 Sout<0> 50 64 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.84781e-13 AS=2.30344e-13 PD=1.77e-06 PS=2.04e-06 $X=23315 $Y=2565 $D=0
M111 Sout<2> 51 65 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.84781e-13 AS=2.30344e-13 PD=1.77e-06 PS=2.04e-06 $X=23315 $Y=9965 $D=0
M112 66 44 Sout<0> vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.17687e-13 AS=1.84781e-13 PD=1.965e-06 PS=1.77e-06 $X=24510 $Y=2565 $D=0
M113 67 45 Sout<2> vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.17687e-13 AS=1.84781e-13 PD=1.965e-06 PS=1.77e-06 $X=24510 $Y=9965 $D=0
M114 vdd! C_in 66 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.3625e-13 AS=2.17687e-13 PD=2.075e-06 PS=1.965e-06 $X=25900 $Y=2565 $D=0
M115 vdd! 10 67 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.3625e-13 AS=2.17687e-13 PD=2.075e-06 PS=1.965e-06 $X=25900 $Y=9965 $D=0
M116 vdd! 17 46 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.94062e-13 AS=1.94062e-13 PD=1.825e-06 PS=1.825e-06 $X=26450 $Y=4425 $D=0
M117 vdd! 18 47 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.94062e-13 AS=1.94062e-13 PD=1.825e-06 PS=1.825e-06 $X=26450 $Y=11825 $D=0
M118 vdd! B<1> 48 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.94062e-13 AS=1.94062e-13 PD=1.825e-06 PS=1.825e-06 $X=30335 $Y=4420 $D=0
M119 vdd! B<3> 49 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.94062e-13 AS=1.94062e-13 PD=1.825e-06 PS=1.825e-06 $X=30335 $Y=11820 $D=0
M120 50 C_in vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.94062e-13 AS=1.94062e-13 PD=1.825e-06 PS=1.825e-06 $X=31065 $Y=2635 $D=0
M121 51 10 vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.94062e-13 AS=1.94062e-13 PD=1.825e-06 PS=1.825e-06 $X=31065 $Y=10035 $D=0
M122 52 13 vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.65375e-13 AS=1.34156e-13 PD=1.655e-06 PS=1.47e-06 $X=34290 $Y=2565 $D=0
M123 53 14 vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.65375e-13 AS=1.34156e-13 PD=1.655e-06 PS=1.47e-06 $X=34290 $Y=9965 $D=0
M124 vdd! C_in 52 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.51031e-13 AS=1.65375e-13 PD=1.57e-06 PS=1.655e-06 $X=35370 $Y=2565 $D=0
M125 vdd! 10 53 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.51031e-13 AS=1.65375e-13 PD=1.57e-06 PS=1.655e-06 $X=35370 $Y=9965 $D=0
M126 68 B<1> vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.17687e-13 AS=2.3625e-13 PD=1.965e-06 PS=2.075e-06 $X=35500 $Y=4490 $D=0
M127 69 B<3> vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.17687e-13 AS=2.3625e-13 PD=1.965e-06 PS=2.075e-06 $X=35500 $Y=11890 $D=0
M128 17 54 68 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.84781e-13 AS=2.17687e-13 PD=1.77e-06 PS=1.965e-06 $X=36890 $Y=4490 $D=0
M129 18 55 69 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.84781e-13 AS=2.17687e-13 PD=1.77e-06 PS=1.965e-06 $X=36890 $Y=11890 $D=0
M130 70 48 17 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.30344e-13 AS=1.84781e-13 PD=2.04e-06 PS=1.77e-06 $X=38085 $Y=4490 $D=0
M131 71 49 18 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.30344e-13 AS=1.84781e-13 PD=2.04e-06 PS=1.77e-06 $X=38085 $Y=11890 $D=0
M132 15 52 vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.65375e-13 AS=1.34156e-13 PD=1.655e-06 PS=1.47e-06 $X=38290 $Y=2565 $D=0
M133 16 53 vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.65375e-13 AS=1.34156e-13 PD=1.655e-06 PS=1.47e-06 $X=38290 $Y=9965 $D=0
M134 vdd! 32 15 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.51031e-13 AS=1.65375e-13 PD=1.57e-06 PS=1.655e-06 $X=39370 $Y=2565 $D=0
M135 vdd! 33 16 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.51031e-13 AS=1.65375e-13 PD=1.57e-06 PS=1.655e-06 $X=39370 $Y=9965 $D=0
M136 vdd! A<1> 70 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=7.59375e-14 AS=2.30344e-13 PD=1.125e-06 PS=2.04e-06 $X=39550 $Y=4490 $D=0
M137 vdd! A<3> 71 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=7.59375e-14 AS=2.30344e-13 PD=1.125e-06 PS=2.04e-06 $X=39550 $Y=11890 $D=0
M138 32 A<0> vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.65375e-13 AS=1.34156e-13 PD=1.655e-06 PS=1.47e-06 $X=42290 $Y=2565 $D=0
M139 33 A<2> vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.65375e-13 AS=1.34156e-13 PD=1.655e-06 PS=1.47e-06 $X=42290 $Y=9965 $D=0
M140 vdd! A<1> 54 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.94062e-13 AS=1.94062e-13 PD=1.825e-06 PS=1.825e-06 $X=42950 $Y=4425 $D=0
M141 vdd! A<3> 55 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.94062e-13 AS=1.94062e-13 PD=1.825e-06 PS=1.825e-06 $X=42950 $Y=11825 $D=0
M142 vdd! B<0> 32 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.51031e-13 AS=1.65375e-13 PD=1.57e-06 PS=1.655e-06 $X=43370 $Y=2565 $D=0
M143 vdd! B<2> 33 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.51031e-13 AS=1.65375e-13 PD=1.57e-06 PS=1.655e-06 $X=43370 $Y=9965 $D=0
.ENDS
***************************************

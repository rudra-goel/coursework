* SPICE NETLIST
***************************************

.SUBCKT full_adder_1_bit
** N=0 EP=0 IP=0 FDC=0
.ENDS
***************************************

* SPICE NETLIST
***************************************

.SUBCKT XOR2 A Out B vdd! gnd!
** N=11 EP=5 IP=0 FDC=12
M0 4 A gnd! gnd! NMOS_VTL L=5e-08 W=9e-08 AD=5.175e-14 AS=5.175e-14 PD=1.33e-06 PS=1.33e-06 $X=2050 $Y=790 $D=1
M1 gnd! A 2 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.2285e-13 AS=4.05e-14 PD=1.725e-06 PS=8.1e-07 $X=5450 $Y=900 $D=1
M2 11 8 gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=9.855e-14 AS=1.2285e-13 PD=1.455e-06 PS=1.725e-06 $X=6915 $Y=900 $D=1
M3 Out 4 11 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.161e-13 AS=9.855e-14 PD=1.65e-06 PS=1.455e-06 $X=8110 $Y=900 $D=1
M4 2 B Out gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.26e-13 AS=1.161e-13 PD=1.76e-06 PS=1.65e-06 $X=9500 $Y=900 $D=1
M5 8 B gnd! gnd! NMOS_VTL L=5e-08 W=9e-08 AD=5.175e-14 AS=5.175e-14 PD=1.33e-06 PS=1.33e-06 $X=14665 $Y=795 $D=1
M6 4 A vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.94062e-13 AS=1.94062e-13 PD=1.825e-06 PS=1.825e-06 $X=2050 $Y=2630 $D=0
M7 9 A vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.30344e-13 AS=7.59375e-14 PD=2.04e-06 PS=1.125e-06 $X=5450 $Y=2565 $D=0
M8 Out 8 9 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.84781e-13 AS=2.30344e-13 PD=1.77e-06 PS=2.04e-06 $X=6915 $Y=2565 $D=0
M9 10 4 Out vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.17687e-13 AS=1.84781e-13 PD=1.965e-06 PS=1.77e-06 $X=8110 $Y=2565 $D=0
M10 vdd! B 10 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.3625e-13 AS=2.17687e-13 PD=2.075e-06 PS=1.965e-06 $X=9500 $Y=2565 $D=0
M11 8 B vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.94062e-13 AS=1.94062e-13 PD=1.825e-06 PS=1.825e-06 $X=14665 $Y=2635 $D=0
.ENDS
***************************************

* SPICE NETLIST
***************************************

.SUBCKT full_adder_1_bit A B S C_in C_out gnd! vdd!
** N=25 EP=7 IP=0 FDC=36
M0 9 A gnd! gnd! NMOS_VTL L=5e-08 W=9e-08 AD=5.175e-14 AS=5.175e-14 PD=1.33e-06 PS=1.33e-06 $X=1950 $Y=790 $D=1
M1 gnd! A 2 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.2285e-13 AS=4.05e-14 PD=1.725e-06 PS=8.1e-07 $X=5350 $Y=900 $D=1
M2 21 10 gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=9.855e-14 AS=1.2285e-13 PD=1.455e-06 PS=1.725e-06 $X=6815 $Y=900 $D=1
M3 3 9 21 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.161e-13 AS=9.855e-14 PD=1.65e-06 PS=1.455e-06 $X=8010 $Y=900 $D=1
M4 2 B 3 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.26e-13 AS=1.161e-13 PD=1.76e-06 PS=1.65e-06 $X=9400 $Y=900 $D=1
M5 10 B gnd! gnd! NMOS_VTL L=5e-08 W=9e-08 AD=5.175e-14 AS=5.175e-14 PD=1.33e-06 PS=1.33e-06 $X=14565 $Y=795 $D=1
M6 11 3 gnd! gnd! NMOS_VTL L=5e-08 W=9e-08 AD=5.175e-14 AS=5.175e-14 PD=1.33e-06 PS=1.33e-06 $X=18450 $Y=790 $D=1
M7 gnd! 3 5 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.2285e-13 AS=4.05e-14 PD=1.725e-06 PS=8.1e-07 $X=21850 $Y=900 $D=1
M8 22 12 gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=9.855e-14 AS=1.2285e-13 PD=1.455e-06 PS=1.725e-06 $X=23315 $Y=900 $D=1
M9 S 11 22 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.161e-13 AS=9.855e-14 PD=1.65e-06 PS=1.455e-06 $X=24510 $Y=900 $D=1
M10 5 C_in S gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.26e-13 AS=1.161e-13 PD=1.76e-06 PS=1.65e-06 $X=25900 $Y=900 $D=1
M11 12 C_in gnd! gnd! NMOS_VTL L=5e-08 W=9e-08 AD=5.175e-14 AS=5.175e-14 PD=1.33e-06 PS=1.33e-06 $X=31065 $Y=795 $D=1
M12 23 3 gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=8.82e-14 AS=7.155e-14 PD=1.34e-06 PS=1.155e-06 $X=34290 $Y=695 $D=1
M13 13 C_in 23 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=8.595e-14 AS=8.82e-14 PD=1.315e-06 PS=1.34e-06 $X=35370 $Y=695 $D=1
M14 24 13 gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=8.82e-14 AS=7.155e-14 PD=1.34e-06 PS=1.155e-06 $X=38290 $Y=695 $D=1
M15 C_out 8 24 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=8.595e-14 AS=8.82e-14 PD=1.315e-06 PS=1.34e-06 $X=39370 $Y=695 $D=1
M16 25 A gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=8.82e-14 AS=7.155e-14 PD=1.34e-06 PS=1.155e-06 $X=42290 $Y=695 $D=1
M17 8 B 25 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=8.595e-14 AS=8.82e-14 PD=1.315e-06 PS=1.34e-06 $X=43370 $Y=695 $D=1
M18 9 A vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.94062e-13 AS=1.94062e-13 PD=1.825e-06 PS=1.825e-06 $X=1950 $Y=2630 $D=0
M19 17 A vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.30344e-13 AS=7.59375e-14 PD=2.04e-06 PS=1.125e-06 $X=5350 $Y=2565 $D=0
M20 3 10 17 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.84781e-13 AS=2.30344e-13 PD=1.77e-06 PS=2.04e-06 $X=6815 $Y=2565 $D=0
M21 18 9 3 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.17687e-13 AS=1.84781e-13 PD=1.965e-06 PS=1.77e-06 $X=8010 $Y=2565 $D=0
M22 vdd! B 18 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.3625e-13 AS=2.17687e-13 PD=2.075e-06 PS=1.965e-06 $X=9400 $Y=2565 $D=0
M23 10 B vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.94062e-13 AS=1.94062e-13 PD=1.825e-06 PS=1.825e-06 $X=14565 $Y=2635 $D=0
M24 11 3 vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.94062e-13 AS=1.94062e-13 PD=1.825e-06 PS=1.825e-06 $X=18450 $Y=2630 $D=0
M25 19 3 vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.30344e-13 AS=7.59375e-14 PD=2.04e-06 PS=1.125e-06 $X=21850 $Y=2565 $D=0
M26 S 12 19 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.84781e-13 AS=2.30344e-13 PD=1.77e-06 PS=2.04e-06 $X=23315 $Y=2565 $D=0
M27 20 11 S vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.17687e-13 AS=1.84781e-13 PD=1.965e-06 PS=1.77e-06 $X=24510 $Y=2565 $D=0
M28 vdd! C_in 20 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=2.3625e-13 AS=2.17687e-13 PD=2.075e-06 PS=1.965e-06 $X=25900 $Y=2565 $D=0
M29 12 C_in vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.94062e-13 AS=1.94062e-13 PD=1.825e-06 PS=1.825e-06 $X=31065 $Y=2635 $D=0
M30 13 3 vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.65375e-13 AS=1.34156e-13 PD=1.655e-06 PS=1.47e-06 $X=34290 $Y=2565 $D=0
M31 vdd! C_in 13 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.51031e-13 AS=1.65375e-13 PD=1.57e-06 PS=1.655e-06 $X=35370 $Y=2565 $D=0
M32 C_out 13 vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.65375e-13 AS=1.34156e-13 PD=1.655e-06 PS=1.47e-06 $X=38290 $Y=2565 $D=0
M33 vdd! 8 C_out vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.51031e-13 AS=1.65375e-13 PD=1.57e-06 PS=1.655e-06 $X=39370 $Y=2565 $D=0
M34 8 A vdd! vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.65375e-13 AS=1.34156e-13 PD=1.655e-06 PS=1.47e-06 $X=42290 $Y=2565 $D=0
M35 vdd! B 8 vdd! PMOS_VTL L=5e-08 W=3.375e-07 AD=1.51031e-13 AS=1.65375e-13 PD=1.57e-06 PS=1.655e-06 $X=43370 $Y=2565 $D=0
.ENDS
***************************************
